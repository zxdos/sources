-- ZPU
--
-- Copyright 2004-2008 oharboe - �yvind Harboe - oyvind.harboe@zylin.com
-- Modified by Alastair M. Robinson for the ZPUFlex project.
--
-- The FreeBSD license
-- 
-- Redistribution and use in source and binary forms, with or without
-- modification, are permitted provided that the following conditions
-- are met:
-- 
-- 1. Redistributions of source code must retain the above copyright
--    notice, this list of conditions and the following disclaimer.
-- 2. Redistributions in binary form must reproduce the above
--    copyright notice, this list of conditions and the following
--    disclaimer in the documentation and/or other materials
--    provided with the distribution.
-- 
-- THIS SOFTWARE IS PROVIDED BY THE ZPU PROJECT ``AS IS'' AND ANY
-- EXPRESS OR IMPLIED WARRANTIES, INCLUDING, BUT NOT LIMITED TO,
-- THE IMPLIED WARRANTIES OF MERCHANTABILITY AND FITNESS FOR A
-- PARTICULAR PURPOSE ARE DISCLAIMED. IN NO EVENT SHALL THE
-- ZPU PROJECT OR CONTRIBUTORS BE LIABLE FOR ANY DIRECT,
-- INDIRECT, INCIDENTAL, SPECIAL, EXEMPLARY, OR CONSEQUENTIAL DAMAGES
-- (INCLUDING, BUT NOT LIMITED TO, PROCUREMENT OF SUBSTITUTE GOODS
-- OR SERVICES; LOSS OF USE, DATA, OR PROFITS; OR BUSINESS INTERRUPTION)
-- HOWEVER CAUSED AND ON ANY THEORY OF LIABILITY, WHETHER IN CONTRACT,
-- STRICT LIABILITY, OR TORT (INCLUDING NEGLIGENCE OR OTHERWISE)
-- ARISING IN ANY WAY OUT OF THE USE OF THIS SOFTWARE, EVEN IF
-- ADVISED OF THE POSSIBILITY OF SUCH DAMAGE.
-- 
-- The views and conclusions contained in the software and documentation
-- are those of the authors and should not be interpreted as representing
-- official policies, either expressed or implied, of the ZPU Project.

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;


library work;
use work.zpupkg.all;

entity CtrlROM_ROM is
generic
	(
		maxAddrBitBRAM : integer := maxAddrBitBRAMLimit -- Specify your actual ROM size to save LEs and unnecessary block RAM usage.
	);
port (
	clk : in std_logic;
	areset : in std_logic := '0';
	from_zpu : in ZPU_ToROM;
	to_zpu : out ZPU_FromROM
);
end CtrlROM_ROM;

architecture arch of CtrlROM_ROM is

type ram_type is array(natural range 0 to ((2**(maxAddrBitBRAM+1))/4)-1) of std_logic_vector(wordSize-1 downto 0);

shared variable ram : ram_type :=
(
     0 => x"0b0b0b0b",
     1 => x"8c0b0b0b",
     2 => x"0b81e004",
     3 => x"0b0b0b0b",
     4 => x"8c04ff0d",
     5 => x"80040400",
     6 => x"00000016",
     7 => x"00000000",
     8 => x"0b0b0bab",
     9 => x"d0080b0b",
    10 => x"0babd408",
    11 => x"0b0b0bab",
    12 => x"d8080b0b",
    13 => x"0b0b9808",
    14 => x"2d0b0b0b",
    15 => x"abd80c0b",
    16 => x"0b0babd4",
    17 => x"0c0b0b0b",
    18 => x"abd00c04",
    19 => x"00000000",
    20 => x"00000000",
    21 => x"00000000",
    22 => x"00000000",
    23 => x"00000000",
    24 => x"71fd0608",
    25 => x"72830609",
    26 => x"81058205",
    27 => x"832b2a83",
    28 => x"ffff0652",
    29 => x"0471fc06",
    30 => x"08728306",
    31 => x"09810583",
    32 => x"05101010",
    33 => x"2a81ff06",
    34 => x"520471fd",
    35 => x"060883ff",
    36 => x"ff738306",
    37 => x"09810582",
    38 => x"05832b2b",
    39 => x"09067383",
    40 => x"ffff0673",
    41 => x"83060981",
    42 => x"05820583",
    43 => x"2b0b2b07",
    44 => x"72fc060c",
    45 => x"51510471",
    46 => x"fc06080b",
    47 => x"0b0ba5ec",
    48 => x"73830610",
    49 => x"10050806",
    50 => x"7381ff06",
    51 => x"73830609",
    52 => x"81058305",
    53 => x"1010102b",
    54 => x"0772fc06",
    55 => x"0c515104",
    56 => x"abd070b0",
    57 => x"ec278b38",
    58 => x"80717084",
    59 => x"05530c81",
    60 => x"e2048c51",
    61 => x"85e80402",
    62 => x"fc050df8",
    63 => x"80518f0b",
    64 => x"abe00c9f",
    65 => x"0babe40c",
    66 => x"a0717081",
    67 => x"055334ab",
    68 => x"e408ff05",
    69 => x"abe40cab",
    70 => x"e4088025",
    71 => x"eb38abe0",
    72 => x"08ff05ab",
    73 => x"e00cabe0",
    74 => x"088025d7",
    75 => x"38800bab",
    76 => x"e40c800b",
    77 => x"abe00c02",
    78 => x"84050d04",
    79 => x"02f0050d",
    80 => x"f88053f8",
    81 => x"a05483bf",
    82 => x"52737081",
    83 => x"05553351",
    84 => x"70737081",
    85 => x"055534ff",
    86 => x"12527180",
    87 => x"25eb38fb",
    88 => x"c0539f52",
    89 => x"a0737081",
    90 => x"055534ff",
    91 => x"12527180",
    92 => x"25f23802",
    93 => x"90050d04",
    94 => x"02f4050d",
    95 => x"74538e0b",
    96 => x"abe00825",
    97 => x"8f3882bc",
    98 => x"2dabe008",
    99 => x"ff05abe0",
   100 => x"0c82fe04",
   101 => x"abe008ab",
   102 => x"e4085351",
   103 => x"728a2e09",
   104 => x"8106b738",
   105 => x"7151719f",
   106 => x"24a038ab",
   107 => x"e008a029",
   108 => x"11f88011",
   109 => x"5151a071",
   110 => x"34abe408",
   111 => x"8105abe4",
   112 => x"0cabe408",
   113 => x"519f7125",
   114 => x"e238800b",
   115 => x"abe40cab",
   116 => x"e0088105",
   117 => x"abe00c83",
   118 => x"ee0470a0",
   119 => x"2912f880",
   120 => x"11515172",
   121 => x"7134abe4",
   122 => x"088105ab",
   123 => x"e40cabe4",
   124 => x"08a02e09",
   125 => x"81068e38",
   126 => x"800babe4",
   127 => x"0cabe008",
   128 => x"8105abe0",
   129 => x"0c028c05",
   130 => x"0d0402ec",
   131 => x"050d800b",
   132 => x"abe80cf6",
   133 => x"8c08f690",
   134 => x"0871882c",
   135 => x"565481ff",
   136 => x"06527372",
   137 => x"25883871",
   138 => x"54820bab",
   139 => x"e80c7288",
   140 => x"2c7381ff",
   141 => x"06545574",
   142 => x"73258b38",
   143 => x"72abe808",
   144 => x"8407abe8",
   145 => x"0c557384",
   146 => x"2b86a071",
   147 => x"25837131",
   148 => x"700b0b0b",
   149 => x"a9a40c81",
   150 => x"712bff05",
   151 => x"f6880cfc",
   152 => x"08fe9014",
   153 => x"ff132c79",
   154 => x"8829fed0",
   155 => x"0570812c",
   156 => x"abe80852",
   157 => x"59535155",
   158 => x"51525476",
   159 => x"802e8538",
   160 => x"70810751",
   161 => x"70f6940c",
   162 => x"71098105",
   163 => x"f6800c72",
   164 => x"098105f6",
   165 => x"840c0294",
   166 => x"050d0402",
   167 => x"f4050d74",
   168 => x"53727081",
   169 => x"055480f5",
   170 => x"2d527180",
   171 => x"2e893871",
   172 => x"5182f82d",
   173 => x"85a10481",
   174 => x"0babd00c",
   175 => x"028c050d",
   176 => x"0402fc05",
   177 => x"0d818080",
   178 => x"51c01151",
   179 => x"70fb3802",
   180 => x"84050d04",
   181 => x"02fc050d",
   182 => x"ec518371",
   183 => x"0c85c12d",
   184 => x"82710c02",
   185 => x"84050d04",
   186 => x"02f0050d",
   187 => x"805185d4",
   188 => x"2d840bec",
   189 => x"0c8ba02d",
   190 => x"87e72d81",
   191 => x"f72d8352",
   192 => x"8b852d81",
   193 => x"51848a2d",
   194 => x"ff125271",
   195 => x"8025f138",
   196 => x"840bec0c",
   197 => x"a7e05185",
   198 => x"9b2d9fdd",
   199 => x"2dabd008",
   200 => x"802e81ae",
   201 => x"38bf0bab",
   202 => x"a00cbf0b",
   203 => x"fc0ca9a8",
   204 => x"518deb2d",
   205 => x"8bcf2d87",
   206 => x"f32d8dfb",
   207 => x"2daa900b",
   208 => x"80f52d70",
   209 => x"872baba0",
   210 => x"08708106",
   211 => x"53565452",
   212 => x"71802e85",
   213 => x"38728107",
   214 => x"5373812a",
   215 => x"70810651",
   216 => x"5271802e",
   217 => x"85387282",
   218 => x"07537382",
   219 => x"2a708106",
   220 => x"51527180",
   221 => x"2e853872",
   222 => x"84075373",
   223 => x"832a7081",
   224 => x"06515271",
   225 => x"802e8538",
   226 => x"72880753",
   227 => x"73842a70",
   228 => x"81065152",
   229 => x"71802e85",
   230 => x"38729007",
   231 => x"5373852a",
   232 => x"70810651",
   233 => x"5271802e",
   234 => x"853872a0",
   235 => x"07537386",
   236 => x"2a708106",
   237 => x"51527180",
   238 => x"2e863872",
   239 => x"80c00753",
   240 => x"72fc0c86",
   241 => x"52abd008",
   242 => x"83388452",
   243 => x"71ec0c86",
   244 => x"b704800b",
   245 => x"abd00c02",
   246 => x"90050d04",
   247 => x"71980c04",
   248 => x"ffb008ab",
   249 => x"d00c0481",
   250 => x"0bffb00c",
   251 => x"04800bff",
   252 => x"b00c0402",
   253 => x"f4050d88",
   254 => x"f504abd0",
   255 => x"0881f02e",
   256 => x"09810689",
   257 => x"38810bab",
   258 => x"980c88f5",
   259 => x"04abd008",
   260 => x"81e02e09",
   261 => x"81068938",
   262 => x"810bab9c",
   263 => x"0c88f504",
   264 => x"abd00852",
   265 => x"ab9c0880",
   266 => x"2e8838ab",
   267 => x"d0088180",
   268 => x"05527184",
   269 => x"2c728f06",
   270 => x"5353ab98",
   271 => x"08802e99",
   272 => x"38728429",
   273 => x"aad80572",
   274 => x"1381712b",
   275 => x"70097308",
   276 => x"06730c51",
   277 => x"535388eb",
   278 => x"04728429",
   279 => x"aad80572",
   280 => x"1383712b",
   281 => x"72080772",
   282 => x"0c535380",
   283 => x"0bab9c0c",
   284 => x"800bab98",
   285 => x"0cabec51",
   286 => x"89f62dab",
   287 => x"d008ff24",
   288 => x"fef83880",
   289 => x"0babd00c",
   290 => x"028c050d",
   291 => x"0402f805",
   292 => x"0daad852",
   293 => x"8f518072",
   294 => x"70840554",
   295 => x"0cff1151",
   296 => x"708025f2",
   297 => x"38028805",
   298 => x"0d0402f0",
   299 => x"050d7551",
   300 => x"87ed2d70",
   301 => x"822cfc06",
   302 => x"aad81172",
   303 => x"109e0671",
   304 => x"0870722a",
   305 => x"70830682",
   306 => x"742b7009",
   307 => x"7406760c",
   308 => x"54515657",
   309 => x"53515387",
   310 => x"e72d71ab",
   311 => x"d00c0290",
   312 => x"050d0402",
   313 => x"fc050d72",
   314 => x"5180710c",
   315 => x"800b8412",
   316 => x"0c028405",
   317 => x"0d0402f0",
   318 => x"050d7570",
   319 => x"08841208",
   320 => x"535353ff",
   321 => x"5471712e",
   322 => x"a83887ed",
   323 => x"2d841308",
   324 => x"70842914",
   325 => x"88117008",
   326 => x"7081ff06",
   327 => x"84180881",
   328 => x"11870684",
   329 => x"1a0c5351",
   330 => x"55515151",
   331 => x"87e72d71",
   332 => x"5473abd0",
   333 => x"0c029005",
   334 => x"0d0402f4",
   335 => x"050d87ed",
   336 => x"2de00870",
   337 => x"8b2a7081",
   338 => x"06515253",
   339 => x"70802e9d",
   340 => x"38abec08",
   341 => x"708429ab",
   342 => x"f4057481",
   343 => x"ff06710c",
   344 => x"5151abec",
   345 => x"08811187",
   346 => x"06abec0c",
   347 => x"51728c2c",
   348 => x"bf06ac94",
   349 => x"0c800bac",
   350 => x"980c87e0",
   351 => x"2d87e72d",
   352 => x"028c050d",
   353 => x"0402fc05",
   354 => x"0d87ed2d",
   355 => x"810bac98",
   356 => x"0c87e72d",
   357 => x"ac980851",
   358 => x"70fa3802",
   359 => x"84050d04",
   360 => x"02fc050d",
   361 => x"abec5189",
   362 => x"e32d898d",
   363 => x"2d8aba51",
   364 => x"87dc2d02",
   365 => x"84050d04",
   366 => x"02fc050d",
   367 => x"8fcf5185",
   368 => x"c12dff11",
   369 => x"51708025",
   370 => x"f6380284",
   371 => x"050d0402",
   372 => x"fc050d81",
   373 => x"0babcc0c",
   374 => x"8151848a",
   375 => x"2d028405",
   376 => x"0d0402fc",
   377 => x"050d8bec",
   378 => x"0487f32d",
   379 => x"80f65189",
   380 => x"aa2dabd0",
   381 => x"08f33880",
   382 => x"da5189aa",
   383 => x"2dabd008",
   384 => x"e838abc8",
   385 => x"085189aa",
   386 => x"2dabd008",
   387 => x"dc38abd0",
   388 => x"08abcc0c",
   389 => x"abd00851",
   390 => x"848a2d02",
   391 => x"84050d04",
   392 => x"02ec050d",
   393 => x"76548052",
   394 => x"870b8815",
   395 => x"80f52d56",
   396 => x"53747224",
   397 => x"8338a053",
   398 => x"725182f8",
   399 => x"2d81128b",
   400 => x"1580f52d",
   401 => x"54527272",
   402 => x"25de3802",
   403 => x"94050d04",
   404 => x"02f0050d",
   405 => x"aca00854",
   406 => x"81f72d80",
   407 => x"0baca40c",
   408 => x"7308802e",
   409 => x"81803882",
   410 => x"0babe40c",
   411 => x"aca4088f",
   412 => x"06abe00c",
   413 => x"73085271",
   414 => x"832e9638",
   415 => x"71832689",
   416 => x"3871812e",
   417 => x"af388dd1",
   418 => x"0471852e",
   419 => x"9f388dd1",
   420 => x"04881480",
   421 => x"f52d8415",
   422 => x"08a7f853",
   423 => x"5452859b",
   424 => x"2d718429",
   425 => x"13700852",
   426 => x"528dd504",
   427 => x"73518ca0",
   428 => x"2d8dd104",
   429 => x"aba00888",
   430 => x"15082c70",
   431 => x"81065152",
   432 => x"71802e87",
   433 => x"38a7fc51",
   434 => x"8dce04a8",
   435 => x"8051859b",
   436 => x"2d841408",
   437 => x"51859b2d",
   438 => x"aca40881",
   439 => x"05aca40c",
   440 => x"8c14548c",
   441 => x"e0040290",
   442 => x"050d0471",
   443 => x"aca00c8c",
   444 => x"d02daca4",
   445 => x"08ff05ac",
   446 => x"a80c0402",
   447 => x"e8050dac",
   448 => x"a008acac",
   449 => x"08575580",
   450 => x"f65189aa",
   451 => x"2dabd008",
   452 => x"812a7081",
   453 => x"06515271",
   454 => x"802e9f38",
   455 => x"8ea20487",
   456 => x"f32d80f6",
   457 => x"5189aa2d",
   458 => x"abd008f3",
   459 => x"38abcc08",
   460 => x"813270ab",
   461 => x"cc0c5184",
   462 => x"8a2d800b",
   463 => x"ac9c0c8c",
   464 => x"5189aa2d",
   465 => x"abd00881",
   466 => x"2a708106",
   467 => x"51527180",
   468 => x"2ebd38ab",
   469 => x"a408abb8",
   470 => x"08aba40c",
   471 => x"abb80cab",
   472 => x"a808abbc",
   473 => x"08aba80c",
   474 => x"abbc0cab",
   475 => x"ac08abc0",
   476 => x"08abac0c",
   477 => x"abc00cab",
   478 => x"b008abc4",
   479 => x"08abb00c",
   480 => x"abc40cab",
   481 => x"b408abc8",
   482 => x"08abb40c",
   483 => x"abc80cac",
   484 => x"9408a006",
   485 => x"52807225",
   486 => x"96388bb8",
   487 => x"2d87f32d",
   488 => x"abcc0881",
   489 => x"3270abcc",
   490 => x"0c705252",
   491 => x"848a2dab",
   492 => x"cc0881ea",
   493 => x"38abb808",
   494 => x"5189aa2d",
   495 => x"abd00880",
   496 => x"2e8938ac",
   497 => x"9c088107",
   498 => x"ac9c0cab",
   499 => x"bc085189",
   500 => x"aa2dabd0",
   501 => x"08802e89",
   502 => x"38ac9c08",
   503 => x"8207ac9c",
   504 => x"0cabc008",
   505 => x"5189aa2d",
   506 => x"abd00880",
   507 => x"2e8938ac",
   508 => x"9c088407",
   509 => x"ac9c0cab",
   510 => x"c4085189",
   511 => x"aa2dabd0",
   512 => x"08802e89",
   513 => x"38ac9c08",
   514 => x"8807ac9c",
   515 => x"0cabc808",
   516 => x"5189aa2d",
   517 => x"abd00880",
   518 => x"2e8938ac",
   519 => x"9c089007",
   520 => x"ac9c0cab",
   521 => x"a4085189",
   522 => x"aa2dabd0",
   523 => x"08802e8a",
   524 => x"38ac9c08",
   525 => x"828007ac",
   526 => x"9c0caba8",
   527 => x"085189aa",
   528 => x"2dabd008",
   529 => x"802e8a38",
   530 => x"ac9c0884",
   531 => x"8007ac9c",
   532 => x"0cabac08",
   533 => x"5189aa2d",
   534 => x"abd00880",
   535 => x"2e8a38ac",
   536 => x"9c088880",
   537 => x"07ac9c0c",
   538 => x"abb00851",
   539 => x"89aa2dab",
   540 => x"d008802e",
   541 => x"8a38ac9c",
   542 => x"08908007",
   543 => x"ac9c0cab",
   544 => x"b4085189",
   545 => x"aa2dabd0",
   546 => x"08802e8a",
   547 => x"38ac9c08",
   548 => x"a08007ac",
   549 => x"9c0cac9c",
   550 => x"08ed0c97",
   551 => x"e40481f5",
   552 => x"5189aa2d",
   553 => x"abd00881",
   554 => x"2a708106",
   555 => x"515271a0",
   556 => x"38abb808",
   557 => x"5189aa2d",
   558 => x"abd00881",
   559 => x"2a708106",
   560 => x"5152718c",
   561 => x"38ac9408",
   562 => x"90065280",
   563 => x"7225bd38",
   564 => x"ac940890",
   565 => x"06528072",
   566 => x"2584388b",
   567 => x"b82daca8",
   568 => x"08527180",
   569 => x"2e8938ff",
   570 => x"12aca80c",
   571 => x"928c04ac",
   572 => x"a40810ac",
   573 => x"a4080570",
   574 => x"84291651",
   575 => x"52881208",
   576 => x"802e8938",
   577 => x"ff518812",
   578 => x"0852712d",
   579 => x"81f25189",
   580 => x"aa2dabd0",
   581 => x"08812a70",
   582 => x"81065152",
   583 => x"71a038ab",
   584 => x"bc085189",
   585 => x"aa2dabd0",
   586 => x"08812a70",
   587 => x"81065152",
   588 => x"718c38ac",
   589 => x"94088806",
   590 => x"52807225",
   591 => x"bf38ac94",
   592 => x"08880652",
   593 => x"80722584",
   594 => x"388bb82d",
   595 => x"aca408ff",
   596 => x"11aca808",
   597 => x"56535373",
   598 => x"72258938",
   599 => x"8114aca8",
   600 => x"0c92fc04",
   601 => x"72101370",
   602 => x"84291651",
   603 => x"52881208",
   604 => x"802e8938",
   605 => x"fe518812",
   606 => x"0852712d",
   607 => x"81fd5189",
   608 => x"aa2dabd0",
   609 => x"08812a70",
   610 => x"81065152",
   611 => x"719738ab",
   612 => x"c0085189",
   613 => x"aa2dabd0",
   614 => x"08812a70",
   615 => x"81065152",
   616 => x"71802ead",
   617 => x"38aca808",
   618 => x"802e8938",
   619 => x"800baca8",
   620 => x"0c93d104",
   621 => x"aca40810",
   622 => x"aca40805",
   623 => x"70842916",
   624 => x"51528812",
   625 => x"08802e89",
   626 => x"38fd5188",
   627 => x"12085271",
   628 => x"2d81fa51",
   629 => x"89aa2dab",
   630 => x"d008812a",
   631 => x"70810651",
   632 => x"52719738",
   633 => x"abc40851",
   634 => x"89aa2dab",
   635 => x"d008812a",
   636 => x"70810651",
   637 => x"5271802e",
   638 => x"ae38aca4",
   639 => x"08ff1154",
   640 => x"52aca808",
   641 => x"73258838",
   642 => x"72aca80c",
   643 => x"94a70471",
   644 => x"10127084",
   645 => x"29165152",
   646 => x"88120880",
   647 => x"2e8938fc",
   648 => x"51881208",
   649 => x"52712dac",
   650 => x"a8087053",
   651 => x"5473802e",
   652 => x"8a388c15",
   653 => x"ff155555",
   654 => x"94ad0482",
   655 => x"0babe40c",
   656 => x"718f06ab",
   657 => x"e00c81eb",
   658 => x"5189aa2d",
   659 => x"abd00881",
   660 => x"2a708106",
   661 => x"51527180",
   662 => x"2ead3874",
   663 => x"08852e09",
   664 => x"8106a438",
   665 => x"881580f5",
   666 => x"2dff0552",
   667 => x"71881681",
   668 => x"b72d7198",
   669 => x"2b527180",
   670 => x"25883880",
   671 => x"0b881681",
   672 => x"b72d7451",
   673 => x"8ca02d81",
   674 => x"f45189aa",
   675 => x"2dabd008",
   676 => x"812a7081",
   677 => x"06515271",
   678 => x"802eb338",
   679 => x"7408852e",
   680 => x"098106aa",
   681 => x"38881580",
   682 => x"f52d8105",
   683 => x"52718816",
   684 => x"81b72d71",
   685 => x"81ff068b",
   686 => x"1680f52d",
   687 => x"54527272",
   688 => x"27873872",
   689 => x"881681b7",
   690 => x"2d74518c",
   691 => x"a02d80da",
   692 => x"5189aa2d",
   693 => x"abd00881",
   694 => x"2a708106",
   695 => x"5152718d",
   696 => x"38ac9408",
   697 => x"81065280",
   698 => x"722581b4",
   699 => x"38aca008",
   700 => x"ac940881",
   701 => x"06535380",
   702 => x"72258438",
   703 => x"8bb82dac",
   704 => x"a8085473",
   705 => x"802e8a38",
   706 => x"8c13ff15",
   707 => x"55539683",
   708 => x"04720852",
   709 => x"71822ea6",
   710 => x"38718226",
   711 => x"89387181",
   712 => x"2ea93897",
   713 => x"a0047183",
   714 => x"2eb13871",
   715 => x"842e0981",
   716 => x"0680ed38",
   717 => x"88130851",
   718 => x"8deb2d97",
   719 => x"a004aca8",
   720 => x"08518813",
   721 => x"0852712d",
   722 => x"97a00481",
   723 => x"0b881408",
   724 => x"2baba008",
   725 => x"32aba00c",
   726 => x"96f60488",
   727 => x"1380f52d",
   728 => x"81058b14",
   729 => x"80f52d53",
   730 => x"54717424",
   731 => x"83388054",
   732 => x"73881481",
   733 => x"b72d8cd0",
   734 => x"2d97a004",
   735 => x"7508802e",
   736 => x"a2387508",
   737 => x"5189aa2d",
   738 => x"abd00881",
   739 => x"06527180",
   740 => x"2e8b38ac",
   741 => x"a8085184",
   742 => x"16085271",
   743 => x"2d881656",
   744 => x"75da3880",
   745 => x"54800bab",
   746 => x"e40c738f",
   747 => x"06abe00c",
   748 => x"a05273ac",
   749 => x"a8082e09",
   750 => x"81069838",
   751 => x"aca408ff",
   752 => x"05743270",
   753 => x"09810570",
   754 => x"72079f2a",
   755 => x"91713151",
   756 => x"51535371",
   757 => x"5182f82d",
   758 => x"8114548e",
   759 => x"7425c638",
   760 => x"abcc0852",
   761 => x"71abd00c",
   762 => x"0298050d",
   763 => x"0402f405",
   764 => x"0dd45281",
   765 => x"ff720c71",
   766 => x"085381ff",
   767 => x"720c7288",
   768 => x"2b83fe80",
   769 => x"06720870",
   770 => x"81ff0651",
   771 => x"525381ff",
   772 => x"720c7271",
   773 => x"07882b72",
   774 => x"087081ff",
   775 => x"06515253",
   776 => x"81ff720c",
   777 => x"72710788",
   778 => x"2b720870",
   779 => x"81ff0672",
   780 => x"07abd00c",
   781 => x"5253028c",
   782 => x"050d0402",
   783 => x"f4050d74",
   784 => x"767181ff",
   785 => x"06d40c53",
   786 => x"53acb008",
   787 => x"85387189",
   788 => x"2b527198",
   789 => x"2ad40c71",
   790 => x"902a7081",
   791 => x"ff06d40c",
   792 => x"5171882a",
   793 => x"7081ff06",
   794 => x"d40c5171",
   795 => x"81ff06d4",
   796 => x"0c72902a",
   797 => x"7081ff06",
   798 => x"d40c51d4",
   799 => x"087081ff",
   800 => x"06515182",
   801 => x"b8bf5270",
   802 => x"81ff2e09",
   803 => x"81069438",
   804 => x"81ff0bd4",
   805 => x"0cd40870",
   806 => x"81ff06ff",
   807 => x"14545151",
   808 => x"71e53870",
   809 => x"abd00c02",
   810 => x"8c050d04",
   811 => x"02fc050d",
   812 => x"81c75181",
   813 => x"ff0bd40c",
   814 => x"ff115170",
   815 => x"8025f438",
   816 => x"0284050d",
   817 => x"0402f405",
   818 => x"0d81ff0b",
   819 => x"d40c9353",
   820 => x"805287fc",
   821 => x"80c15198",
   822 => x"bb2dabd0",
   823 => x"088b3881",
   824 => x"ff0bd40c",
   825 => x"815399f2",
   826 => x"0499ac2d",
   827 => x"ff135372",
   828 => x"df3872ab",
   829 => x"d00c028c",
   830 => x"050d0402",
   831 => x"ec050d81",
   832 => x"0bacb00c",
   833 => x"8454d008",
   834 => x"708f2a70",
   835 => x"81065151",
   836 => x"5372f338",
   837 => x"72d00c99",
   838 => x"ac2da884",
   839 => x"51859b2d",
   840 => x"d008708f",
   841 => x"2a708106",
   842 => x"51515372",
   843 => x"f338810b",
   844 => x"d00cb153",
   845 => x"805284d4",
   846 => x"80c05198",
   847 => x"bb2dabd0",
   848 => x"08812e93",
   849 => x"3872822e",
   850 => x"bd38ff13",
   851 => x"5372e538",
   852 => x"ff145473",
   853 => x"ffb03899",
   854 => x"ac2d83aa",
   855 => x"52849c80",
   856 => x"c85198bb",
   857 => x"2dabd008",
   858 => x"812e0981",
   859 => x"06923897",
   860 => x"ed2dabd0",
   861 => x"0883ffff",
   862 => x"06537283",
   863 => x"aa2e9d38",
   864 => x"99c52d9b",
   865 => x"9704a890",
   866 => x"51859b2d",
   867 => x"80539ce5",
   868 => x"04a8a851",
   869 => x"859b2d80",
   870 => x"549cb704",
   871 => x"81ff0bd4",
   872 => x"0cb15499",
   873 => x"ac2d8fcf",
   874 => x"53805287",
   875 => x"fc80f751",
   876 => x"98bb2dab",
   877 => x"d00855ab",
   878 => x"d008812e",
   879 => x"0981069b",
   880 => x"3881ff0b",
   881 => x"d40c820a",
   882 => x"52849c80",
   883 => x"e95198bb",
   884 => x"2dabd008",
   885 => x"802e8d38",
   886 => x"99ac2dff",
   887 => x"135372c9",
   888 => x"389caa04",
   889 => x"81ff0bd4",
   890 => x"0cabd008",
   891 => x"5287fc80",
   892 => x"fa5198bb",
   893 => x"2dabd008",
   894 => x"b13881ff",
   895 => x"0bd40cd4",
   896 => x"085381ff",
   897 => x"0bd40c81",
   898 => x"ff0bd40c",
   899 => x"81ff0bd4",
   900 => x"0c81ff0b",
   901 => x"d40c7286",
   902 => x"2a708106",
   903 => x"76565153",
   904 => x"729538ab",
   905 => x"d008549c",
   906 => x"b7047382",
   907 => x"2efee238",
   908 => x"ff145473",
   909 => x"feed3873",
   910 => x"acb00c73",
   911 => x"8b388152",
   912 => x"87fc80d0",
   913 => x"5198bb2d",
   914 => x"81ff0bd4",
   915 => x"0cd00870",
   916 => x"8f2a7081",
   917 => x"06515153",
   918 => x"72f33872",
   919 => x"d00c81ff",
   920 => x"0bd40c81",
   921 => x"5372abd0",
   922 => x"0c029405",
   923 => x"0d0402e8",
   924 => x"050d7855",
   925 => x"805681ff",
   926 => x"0bd40cd0",
   927 => x"08708f2a",
   928 => x"70810651",
   929 => x"515372f3",
   930 => x"3882810b",
   931 => x"d00c81ff",
   932 => x"0bd40c77",
   933 => x"5287fc80",
   934 => x"d15198bb",
   935 => x"2d80dbc6",
   936 => x"df54abd0",
   937 => x"08802e8a",
   938 => x"38a8c851",
   939 => x"859b2d9e",
   940 => x"850481ff",
   941 => x"0bd40cd4",
   942 => x"087081ff",
   943 => x"06515372",
   944 => x"81fe2e09",
   945 => x"81069d38",
   946 => x"80ff5397",
   947 => x"ed2dabd0",
   948 => x"08757084",
   949 => x"05570cff",
   950 => x"13537280",
   951 => x"25ed3881",
   952 => x"569dea04",
   953 => x"ff145473",
   954 => x"c93881ff",
   955 => x"0bd40c81",
   956 => x"ff0bd40c",
   957 => x"d008708f",
   958 => x"2a708106",
   959 => x"51515372",
   960 => x"f33872d0",
   961 => x"0c75abd0",
   962 => x"0c029805",
   963 => x"0d0402e8",
   964 => x"050d7779",
   965 => x"7b585555",
   966 => x"80537276",
   967 => x"25a33874",
   968 => x"70810556",
   969 => x"80f52d74",
   970 => x"70810556",
   971 => x"80f52d52",
   972 => x"5271712e",
   973 => x"86388151",
   974 => x"9ec30481",
   975 => x"13539e9a",
   976 => x"04805170",
   977 => x"abd00c02",
   978 => x"98050d04",
   979 => x"02ec050d",
   980 => x"76557480",
   981 => x"2ebb389a",
   982 => x"1580e02d",
   983 => x"51a5d02d",
   984 => x"abd008ab",
   985 => x"d008b0e0",
   986 => x"0cabd008",
   987 => x"5454b0bc",
   988 => x"08802e99",
   989 => x"38941580",
   990 => x"e02d51a5",
   991 => x"d02dabd0",
   992 => x"08902b83",
   993 => x"fff00a06",
   994 => x"70750751",
   995 => x"5372b0e0",
   996 => x"0cb0e008",
   997 => x"5372802e",
   998 => x"9938b0b4",
   999 => x"08fe1471",
  1000 => x"29b0c808",
  1001 => x"05b0e40c",
  1002 => x"70842bb0",
  1003 => x"c00c549f",
  1004 => x"d804b0cc",
  1005 => x"08b0e00c",
  1006 => x"b0d008b0",
  1007 => x"e40cb0bc",
  1008 => x"08802e8a",
  1009 => x"38b0b408",
  1010 => x"842b539f",
  1011 => x"d404b0d4",
  1012 => x"08842b53",
  1013 => x"72b0c00c",
  1014 => x"0294050d",
  1015 => x"0402d805",
  1016 => x"0d800bb0",
  1017 => x"bc0c8454",
  1018 => x"99fb2dab",
  1019 => x"d008802e",
  1020 => x"9538acb4",
  1021 => x"5280519c",
  1022 => x"ee2dabd0",
  1023 => x"08802e86",
  1024 => x"38fe54a0",
  1025 => x"8e04ff14",
  1026 => x"54738024",
  1027 => x"db38738c",
  1028 => x"38a8d851",
  1029 => x"859b2d73",
  1030 => x"55a59704",
  1031 => x"8056810b",
  1032 => x"b0e80c88",
  1033 => x"53a8ec52",
  1034 => x"acea519e",
  1035 => x"8e2dabd0",
  1036 => x"08762e09",
  1037 => x"81068738",
  1038 => x"abd008b0",
  1039 => x"e80c8853",
  1040 => x"a8f852ad",
  1041 => x"86519e8e",
  1042 => x"2dabd008",
  1043 => x"8738abd0",
  1044 => x"08b0e80c",
  1045 => x"b0e80880",
  1046 => x"2e80f638",
  1047 => x"affa0b80",
  1048 => x"f52daffb",
  1049 => x"0b80f52d",
  1050 => x"71982b71",
  1051 => x"902b07af",
  1052 => x"fc0b80f5",
  1053 => x"2d70882b",
  1054 => x"7207affd",
  1055 => x"0b80f52d",
  1056 => x"7107b0b2",
  1057 => x"0b80f52d",
  1058 => x"b0b30b80",
  1059 => x"f52d7188",
  1060 => x"2b07535f",
  1061 => x"54525a56",
  1062 => x"57557381",
  1063 => x"abaa2e09",
  1064 => x"81068d38",
  1065 => x"7551a5a0",
  1066 => x"2dabd008",
  1067 => x"56a1bd04",
  1068 => x"7382d4d5",
  1069 => x"2e8738a9",
  1070 => x"8451a1fe",
  1071 => x"04acb452",
  1072 => x"75519cee",
  1073 => x"2dabd008",
  1074 => x"55abd008",
  1075 => x"802e83c7",
  1076 => x"388853a8",
  1077 => x"f852ad86",
  1078 => x"519e8e2d",
  1079 => x"abd00889",
  1080 => x"38810bb0",
  1081 => x"bc0ca284",
  1082 => x"048853a8",
  1083 => x"ec52acea",
  1084 => x"519e8e2d",
  1085 => x"abd00880",
  1086 => x"2e8a38a9",
  1087 => x"9851859b",
  1088 => x"2da2de04",
  1089 => x"b0b20b80",
  1090 => x"f52d5473",
  1091 => x"80d52e09",
  1092 => x"810680ca",
  1093 => x"38b0b30b",
  1094 => x"80f52d54",
  1095 => x"7381aa2e",
  1096 => x"098106ba",
  1097 => x"38800bac",
  1098 => x"b40b80f5",
  1099 => x"2d565474",
  1100 => x"81e92e83",
  1101 => x"38815474",
  1102 => x"81eb2e8c",
  1103 => x"38805573",
  1104 => x"752e0981",
  1105 => x"0682d038",
  1106 => x"acbf0b80",
  1107 => x"f52d5574",
  1108 => x"8d38acc0",
  1109 => x"0b80f52d",
  1110 => x"5473822e",
  1111 => x"86388055",
  1112 => x"a59704ac",
  1113 => x"c10b80f5",
  1114 => x"2d70b0b4",
  1115 => x"0cff05b0",
  1116 => x"b80cacc2",
  1117 => x"0b80f52d",
  1118 => x"acc30b80",
  1119 => x"f52d5876",
  1120 => x"05778280",
  1121 => x"290570b0",
  1122 => x"c40cacc4",
  1123 => x"0b80f52d",
  1124 => x"70b0d80c",
  1125 => x"b0bc0859",
  1126 => x"57587680",
  1127 => x"2e81a338",
  1128 => x"8853a8f8",
  1129 => x"52ad8651",
  1130 => x"9e8e2dab",
  1131 => x"d00881e7",
  1132 => x"38b0b408",
  1133 => x"70842bb0",
  1134 => x"c00c70b0",
  1135 => x"d40cacd9",
  1136 => x"0b80f52d",
  1137 => x"acd80b80",
  1138 => x"f52d7182",
  1139 => x"802905ac",
  1140 => x"da0b80f5",
  1141 => x"2d708480",
  1142 => x"802912ac",
  1143 => x"db0b80f5",
  1144 => x"2d708180",
  1145 => x"0a291270",
  1146 => x"b0dc0cb0",
  1147 => x"d8087129",
  1148 => x"b0c40805",
  1149 => x"70b0c80c",
  1150 => x"ace10b80",
  1151 => x"f52dace0",
  1152 => x"0b80f52d",
  1153 => x"71828029",
  1154 => x"05ace20b",
  1155 => x"80f52d70",
  1156 => x"84808029",
  1157 => x"12ace30b",
  1158 => x"80f52d70",
  1159 => x"982b81f0",
  1160 => x"0a067205",
  1161 => x"70b0cc0c",
  1162 => x"fe117e29",
  1163 => x"7705b0d0",
  1164 => x"0c525952",
  1165 => x"43545e51",
  1166 => x"5259525d",
  1167 => x"575957a5",
  1168 => x"9004acc6",
  1169 => x"0b80f52d",
  1170 => x"acc50b80",
  1171 => x"f52d7182",
  1172 => x"80290570",
  1173 => x"b0c00c70",
  1174 => x"a02983ff",
  1175 => x"0570892a",
  1176 => x"70b0d40c",
  1177 => x"accb0b80",
  1178 => x"f52dacca",
  1179 => x"0b80f52d",
  1180 => x"71828029",
  1181 => x"0570b0dc",
  1182 => x"0c7b7129",
  1183 => x"1e70b0d0",
  1184 => x"0c7db0cc",
  1185 => x"0c7305b0",
  1186 => x"c80c555e",
  1187 => x"51515555",
  1188 => x"80519ecc",
  1189 => x"2d815574",
  1190 => x"abd00c02",
  1191 => x"a8050d04",
  1192 => x"02f4050d",
  1193 => x"7470882a",
  1194 => x"83fe8006",
  1195 => x"7072982a",
  1196 => x"0772882b",
  1197 => x"87fc8080",
  1198 => x"0673982b",
  1199 => x"81f00a06",
  1200 => x"71730707",
  1201 => x"abd00c56",
  1202 => x"51535102",
  1203 => x"8c050d04",
  1204 => x"02f8050d",
  1205 => x"028e0580",
  1206 => x"f52d7488",
  1207 => x"2b077083",
  1208 => x"ffff06ab",
  1209 => x"d00c5102",
  1210 => x"88050d04",
  1211 => x"00ffffff",
  1212 => x"ff00ffff",
  1213 => x"ffff00ff",
  1214 => x"ffffff00",
  1215 => x"52657365",
  1216 => x"74000000",
  1217 => x"4d616e75",
  1218 => x"616c2053",
  1219 => x"65727665",
  1220 => x"00000000",
  1221 => x"42616c6c",
  1222 => x"20416e67",
  1223 => x"6c650000",
  1224 => x"42616c6c",
  1225 => x"20537065",
  1226 => x"65640000",
  1227 => x"50616464",
  1228 => x"6c652053",
  1229 => x"697a6500",
  1230 => x"536f756e",
  1231 => x"64000000",
  1232 => x"466f7572",
  1233 => x"20706c61",
  1234 => x"79657273",
  1235 => x"00000000",
  1236 => x"446f7562",
  1237 => x"6c65204f",
  1238 => x"53442077",
  1239 => x"696e646f",
  1240 => x"77000000",
  1241 => x"45786974",
  1242 => x"00000000",
  1243 => x"4d6f6e6f",
  1244 => x"00000000",
  1245 => x"47726579",
  1246 => x"7363616c",
  1247 => x"65000000",
  1248 => x"52474231",
  1249 => x"00000000",
  1250 => x"52474232",
  1251 => x"00000000",
  1252 => x"4669656c",
  1253 => x"64000000",
  1254 => x"49636500",
  1255 => x"43687269",
  1256 => x"73746d61",
  1257 => x"73000000",
  1258 => x"4d61726b",
  1259 => x"736d616e",
  1260 => x"00000000",
  1261 => x"4c617320",
  1262 => x"56656761",
  1263 => x"73000000",
  1264 => x"41592d33",
  1265 => x"2d383531",
  1266 => x"3520636f",
  1267 => x"6c6f7273",
  1268 => x"00000000",
  1269 => x"54525120",
  1270 => x"436f6c6f",
  1271 => x"72730000",
  1272 => x"496e6974",
  1273 => x"69616c69",
  1274 => x"7a696e67",
  1275 => x"20534420",
  1276 => x"63617264",
  1277 => x"0a000000",
  1278 => x"16200000",
  1279 => x"14200000",
  1280 => x"15200000",
  1281 => x"53442069",
  1282 => x"6e69742e",
  1283 => x"2e2e0a00",
  1284 => x"53442063",
  1285 => x"61726420",
  1286 => x"72657365",
  1287 => x"74206661",
  1288 => x"696c6564",
  1289 => x"210a0000",
  1290 => x"53444843",
  1291 => x"20657272",
  1292 => x"6f72210a",
  1293 => x"00000000",
  1294 => x"57726974",
  1295 => x"65206661",
  1296 => x"696c6564",
  1297 => x"0a000000",
  1298 => x"52656164",
  1299 => x"20666169",
  1300 => x"6c65640a",
  1301 => x"00000000",
  1302 => x"43617264",
  1303 => x"20696e69",
  1304 => x"74206661",
  1305 => x"696c6564",
  1306 => x"0a000000",
  1307 => x"46415431",
  1308 => x"36202020",
  1309 => x"00000000",
  1310 => x"46415433",
  1311 => x"32202020",
  1312 => x"00000000",
  1313 => x"4e6f2070",
  1314 => x"61727469",
  1315 => x"74696f6e",
  1316 => x"20736967",
  1317 => x"0a000000",
  1318 => x"42616420",
  1319 => x"70617274",
  1320 => x"0a000000",
  1321 => x"00000002",
  1322 => x"00000002",
  1323 => x"000012fc",
  1324 => x"000002d4",
  1325 => x"00000001",
  1326 => x"00001304",
  1327 => x"00000000",
  1328 => x"00000001",
  1329 => x"00001314",
  1330 => x"00000001",
  1331 => x"00000001",
  1332 => x"00001320",
  1333 => x"00000002",
  1334 => x"00000001",
  1335 => x"0000132c",
  1336 => x"00000003",
  1337 => x"00000001",
  1338 => x"00001338",
  1339 => x"00000004",
  1340 => x"00000001",
  1341 => x"00001340",
  1342 => x"00000006",
  1343 => x"00000001",
  1344 => x"00001350",
  1345 => x"00000005",
  1346 => x"00000003",
  1347 => x"0000152c",
  1348 => x"0000000b",
  1349 => x"00000002",
  1350 => x"00001364",
  1351 => x"000005e2",
  1352 => x"00000000",
  1353 => x"00000000",
  1354 => x"00000000",
  1355 => x"0000136c",
  1356 => x"00001374",
  1357 => x"00001380",
  1358 => x"00001388",
  1359 => x"00001390",
  1360 => x"00001398",
  1361 => x"0000139c",
  1362 => x"000013a8",
  1363 => x"000013b4",
  1364 => x"000013c0",
  1365 => x"000013d4",
  1366 => x"00000000",
  1367 => x"00000000",
  1368 => x"00000000",
  1369 => x"00000000",
  1370 => x"00000000",
  1371 => x"00000000",
  1372 => x"00000000",
  1373 => x"00000000",
  1374 => x"00000000",
  1375 => x"00000000",
  1376 => x"00000000",
  1377 => x"00000000",
  1378 => x"00000000",
  1379 => x"00000000",
  1380 => x"00000000",
  1381 => x"00000000",
  1382 => x"00000000",
  1383 => x"00000000",
  1384 => x"00000006",
  1385 => x"00000043",
  1386 => x"00000042",
  1387 => x"0000003b",
  1388 => x"0000004b",
  1389 => x"00000033",
  1390 => x"00000003",
  1391 => x"0000000b",
  1392 => x"00000083",
  1393 => x"00000023",
  1394 => x"0000007e",
  1395 => x"00000000",
	others => x"00000000"
);

begin

process (clk)
begin
	if (clk'event and clk = '1') then
		if (from_zpu.memAWriteEnable = '1') and (from_zpu.memBWriteEnable = '1') and (from_zpu.memAAddr=from_zpu.memBAddr) and (from_zpu.memAWrite/=from_zpu.memBWrite) then
			report "write collision" severity failure;
		end if;
	
		if (from_zpu.memAWriteEnable = '1') then
			ram(to_integer(unsigned(from_zpu.memAAddr(maxAddrBitBRAM downto 2)))) := from_zpu.memAWrite;
			to_zpu.memARead <= from_zpu.memAWrite;
		else
			to_zpu.memARead <= ram(to_integer(unsigned(from_zpu.memAAddr(maxAddrBitBRAM downto 2))));
		end if;
	end if;
end process;

process (clk)
begin
	if (clk'event and clk = '1') then
		if (from_zpu.memBWriteEnable = '1') then
			ram(to_integer(unsigned(from_zpu.memBAddr(maxAddrBitBRAM downto 2)))) := from_zpu.memBWrite;
			to_zpu.memBRead <= from_zpu.memBWrite;
		else
			to_zpu.memBRead <= ram(to_integer(unsigned(from_zpu.memBAddr(maxAddrBitBRAM downto 2))));
		end if;
	end if;
end process;


end arch;

