00
ff
61
2a
62
01
a4
bc
d1
20
61
3a
a4
dc
d1
20
61
4a
a4
fc
d1
20
61
40
62
30
a4
7c
d1
20
61
30
a4
5c
d1
20
62
20
63
30
64
20
6e
01
6d
03
a3
9c
d1
20
a3
bc
61
40
d1
20
65
ff
85
e5
35
00
12
3a
65
ff
85
e5
35
00
12
42
61
30
a3
9c
d1
20
a3
dc
d1
20
65
f0
85
e5
35
00
12
54
d1
20
a3
fc
d1
20
83
d5
84
d5
a4
3c
d3
40
65
f0
85
e5
35
00
12
6a
d3
40
83
d5
84
d5
a4
1c
d3
40
65
f0
85
e5
35
00
12
7c
d3
40
83
d5
84
d5
a4
3c
d3
40
65
f0
85
e5
35
00
12
8e
d3
40
62
00
e2
9e
12
72
00
e0
63
01
61
01
62
07
69
20
6a
0f
65
01
6b
7a
6e
01
6d
00
67
00
a3
98
77
01
47
c0
13
20
62
01
e2
a1
13
10
62
02
e2
a1
13
14
62
04
e2
a1
13
18
62
05
e2
a1
13
1c
62
07
e2
a1
13
74
62
08
e2
a1
13
82
62
0c
e2
a1
13
26
62
0d
e2
a1
13
2c
4c
01
13
74
4c
02
13
82
62
70
82
35
32
00
12
f4
a3
90
c1
3a
6e
40
8e
15
d5
e4
db
e4
4c
01
13
32
4c
02
13
38
12
b4
63
01
12
ea
63
02
12
ea
63
04
12
ea
63
08
12
ea
7d
01
67
00
12
ba
6e
01
8a
e5
12
ea
6e
01
7a
01
12
ea
a3
94
d9
a3
12
b4
a3
98
d9
a3
12
b4
65
08
89
55
8a
55
a5
1c
d9
a0
65
f0
6e
01
85
e5
35
00
13
4c
a5
3c
d9
a0
65
ff
6e
01
85
e5
35
00
13
5a
00
e0
61
2c
62
10
a4
9c
d1
20
61
32
62
25
fd
29
d1
25
12
02
00
fc
a3
94
d9
a3
4f
01
13
3e
6c
01
12
f2
00
fb
a3
98
d9
a3
4f
01
13
3e
6c
02
12
f2
6e
ff
7e
33
e0
7f
e0
00
07
fe
07
99
00
00
20
83
31
86
7f
c7
4a
46
7b
c6
3f
80
5f
43
ff
e4
df
63
ff
e0
db
60
aa
a3
6a
c0
ea
ff
d5
7f
00
00
c6
00
66
00
e6
00
66
00
67
c0
00
00
c0
60
00
84
8c
8e
52
c4
52
84
8c
83
00
00
ff
ff
ff
ff
04
00
1e
03
37
86
7f
87
0f
c6
07
76
0f
f8
0f
db
07
fc
03
ef
01
df
00
9f
00
0f
01
07
ff
ff
ff
7f
00
00
00
03
00
06
00
07
00
06
00
06
00
00
00
03
00
04
00
03
00
00
00
00
00
03
00
00
ff
ff
ff
7f
04
00
1e
00
37
80
7f
80
0f
c0
07
70
0f
f8
0f
d8
07
f8
03
ee
01
df
00
9f
00
4f
00
67
00
03
00
00
10
00
3c
0e
5e
bf
ff
ff
3f
ff
0f
f7
07
fb
07
f9
03
f8
01
fc
00
de
00
9e
00
5f
00
0f
00
0f
00
00
24
30
54
28
54
30
74
29
54
2a
54
29
00
00
50
00
54
80
71
e0
54
80
54
83
54
43
00
00
00
00
00
00
20
02
20
02
20
02
26
c6
aa
aa
26
a6
00
00
70
60
20
a0
24
84
2a
aa
2a
aa
24
64
00
00
00
00
00
00
14
00
14
00
08
94
09
54
08
88
00
00
c4
ee
aa
48
ce
4e
aa
48
aa
48
aa
4e
00
00
07
e0
03
c0
01
80
00
00
ff
7e
ff
7e
e0
18
e0
18
e0
18
fc
18
fc
18
e0
18
e0
18
e0
18
e0
18
e0
7e
e0
7e
00
00
00
00
00
00
ff
70
ff
70
e0
70
e0
70
e0
70
fc
70
fc
70
e0
70
e0
70
e0
70
e0
70
ff
7e
ff
7e
00
00
00
00
00
00
f8
08
fe
1c
e7
3e
e7
3e
e7
3e
e7
3e
e7
1c
e7
1c
e7
1c
e7
08
e7
00
fe
1c
f8
1c
00
00
00
00
00
02
10
0c
08
14
0e
c0
05
a0
06
1c
1a
24
7a
90
c1
e8
02
18
05
08
0c
10
10
00
00
00
00
00
00
00
c3
02
31
8c
09
54
0e
c4
75
b9
1e
1c
1a
3e
7a
93
e1
e9
22
19
05
08
4c
14
30
0a
1b
32
14
32
20
01
