-- ZPU
--
-- Copyright 2004-2008 oharboe - �yvind Harboe - oyvind.harboe@zylin.com
-- Modified by Alastair M. Robinson for the ZPUFlex project.
--
-- The FreeBSD license
-- 
-- Redistribution and use in source and binary forms, with or without
-- modification, are permitted provided that the following conditions
-- are met:
-- 
-- 1. Redistributions of source code must retain the above copyright
--    notice, this list of conditions and the following disclaimer.
-- 2. Redistributions in binary form must reproduce the above
--    copyright notice, this list of conditions and the following
--    disclaimer in the documentation and/or other materials
--    provided with the distribution.
-- 
-- THIS SOFTWARE IS PROVIDED BY THE ZPU PROJECT ``AS IS'' AND ANY
-- EXPRESS OR IMPLIED WARRANTIES, INCLUDING, BUT NOT LIMITED TO,
-- THE IMPLIED WARRANTIES OF MERCHANTABILITY AND FITNESS FOR A
-- PARTICULAR PURPOSE ARE DISCLAIMED. IN NO EVENT SHALL THE
-- ZPU PROJECT OR CONTRIBUTORS BE LIABLE FOR ANY DIRECT,
-- INDIRECT, INCIDENTAL, SPECIAL, EXEMPLARY, OR CONSEQUENTIAL DAMAGES
-- (INCLUDING, BUT NOT LIMITED TO, PROCUREMENT OF SUBSTITUTE GOODS
-- OR SERVICES; LOSS OF USE, DATA, OR PROFITS; OR BUSINESS INTERRUPTION)
-- HOWEVER CAUSED AND ON ANY THEORY OF LIABILITY, WHETHER IN CONTRACT,
-- STRICT LIABILITY, OR TORT (INCLUDING NEGLIGENCE OR OTHERWISE)
-- ARISING IN ANY WAY OUT OF THE USE OF THIS SOFTWARE, EVEN IF
-- ADVISED OF THE POSSIBILITY OF SUCH DAMAGE.
-- 
-- The views and conclusions contained in the software and documentation
-- are those of the authors and should not be interpreted as representing
-- official policies, either expressed or implied, of the ZPU Project.

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;


library work;
use work.zpupkg.all;

entity CtrlROM_ROM is
generic
	(
		maxAddrBitBRAM : integer := maxAddrBitBRAMLimit -- Specify your actual ROM size to save LEs and unnecessary block RAM usage.
	);
port (
	clk : in std_logic;
	areset : in std_logic := '0';
	from_zpu : in ZPU_ToROM;
	to_zpu : out ZPU_FromROM
);
end CtrlROM_ROM;

architecture arch of CtrlROM_ROM is

type ram_type is array(natural range 0 to ((2**(maxAddrBitBRAM+1))/4)-1) of std_logic_vector(wordSize-1 downto 0);

shared variable ram : ram_type :=
(
     0 => x"0b0b0b0b",
     1 => x"8c0b0b0b",
     2 => x"0b81e004",
     3 => x"0b0b0b0b",
     4 => x"8c04ff0d",
     5 => x"80040400",
     6 => x"00000016",
     7 => x"00000000",
     8 => x"0b0b0bae",
     9 => x"f4080b0b",
    10 => x"0baef808",
    11 => x"0b0b0bae",
    12 => x"fc080b0b",
    13 => x"0b0b9808",
    14 => x"2d0b0b0b",
    15 => x"aefc0c0b",
    16 => x"0b0baef8",
    17 => x"0c0b0b0b",
    18 => x"aef40c04",
    19 => x"00000000",
    20 => x"00000000",
    21 => x"00000000",
    22 => x"00000000",
    23 => x"00000000",
    24 => x"71fd0608",
    25 => x"72830609",
    26 => x"81058205",
    27 => x"832b2a83",
    28 => x"ffff0652",
    29 => x"0471fc06",
    30 => x"08728306",
    31 => x"09810583",
    32 => x"05101010",
    33 => x"2a81ff06",
    34 => x"520471fd",
    35 => x"060883ff",
    36 => x"ff738306",
    37 => x"09810582",
    38 => x"05832b2b",
    39 => x"09067383",
    40 => x"ffff0673",
    41 => x"83060981",
    42 => x"05820583",
    43 => x"2b0b2b07",
    44 => x"72fc060c",
    45 => x"51510471",
    46 => x"fc06080b",
    47 => x"0b0ba6c4",
    48 => x"73830610",
    49 => x"10050806",
    50 => x"7381ff06",
    51 => x"73830609",
    52 => x"81058305",
    53 => x"1010102b",
    54 => x"0772fc06",
    55 => x"0c515104",
    56 => x"aef470b4",
    57 => x"90278b38",
    58 => x"80717084",
    59 => x"05530c81",
    60 => x"e2048c51",
    61 => x"85e80402",
    62 => x"fc050df8",
    63 => x"80518f0b",
    64 => x"af840c9f",
    65 => x"0baf880c",
    66 => x"a0717081",
    67 => x"055334af",
    68 => x"8808ff05",
    69 => x"af880caf",
    70 => x"88088025",
    71 => x"eb38af84",
    72 => x"08ff05af",
    73 => x"840caf84",
    74 => x"088025d7",
    75 => x"38800baf",
    76 => x"880c800b",
    77 => x"af840c02",
    78 => x"84050d04",
    79 => x"02f0050d",
    80 => x"f88053f8",
    81 => x"a05483bf",
    82 => x"52737081",
    83 => x"05553351",
    84 => x"70737081",
    85 => x"055534ff",
    86 => x"12527180",
    87 => x"25eb38fb",
    88 => x"c0539f52",
    89 => x"a0737081",
    90 => x"055534ff",
    91 => x"12527180",
    92 => x"25f23802",
    93 => x"90050d04",
    94 => x"02f4050d",
    95 => x"74538e0b",
    96 => x"af840825",
    97 => x"8f3882bc",
    98 => x"2daf8408",
    99 => x"ff05af84",
   100 => x"0c82fe04",
   101 => x"af8408af",
   102 => x"88085351",
   103 => x"728a2e09",
   104 => x"8106b738",
   105 => x"7151719f",
   106 => x"24a038af",
   107 => x"8408a029",
   108 => x"11f88011",
   109 => x"5151a071",
   110 => x"34af8808",
   111 => x"8105af88",
   112 => x"0caf8808",
   113 => x"519f7125",
   114 => x"e238800b",
   115 => x"af880caf",
   116 => x"84088105",
   117 => x"af840c83",
   118 => x"ee0470a0",
   119 => x"2912f880",
   120 => x"11515172",
   121 => x"7134af88",
   122 => x"088105af",
   123 => x"880caf88",
   124 => x"08a02e09",
   125 => x"81068e38",
   126 => x"800baf88",
   127 => x"0caf8408",
   128 => x"8105af84",
   129 => x"0c028c05",
   130 => x"0d0402ec",
   131 => x"050d800b",
   132 => x"af8c0cf6",
   133 => x"8c08f690",
   134 => x"0871882c",
   135 => x"565481ff",
   136 => x"06527372",
   137 => x"25883871",
   138 => x"54820baf",
   139 => x"8c0c7288",
   140 => x"2c7381ff",
   141 => x"06545574",
   142 => x"73258b38",
   143 => x"72af8c08",
   144 => x"8407af8c",
   145 => x"0c557384",
   146 => x"2b86a071",
   147 => x"25827131",
   148 => x"700b0b0b",
   149 => x"ac880c81",
   150 => x"712bff05",
   151 => x"f6880cfc",
   152 => x"08fefe14",
   153 => x"ff132c79",
   154 => x"8829ff94",
   155 => x"0570812c",
   156 => x"af8c0852",
   157 => x"59535155",
   158 => x"51525476",
   159 => x"802e8538",
   160 => x"70810751",
   161 => x"70f6940c",
   162 => x"71098105",
   163 => x"f6800c72",
   164 => x"098105f6",
   165 => x"840c0294",
   166 => x"050d0402",
   167 => x"f4050d74",
   168 => x"53727081",
   169 => x"055480f5",
   170 => x"2d527180",
   171 => x"2e893871",
   172 => x"5182f82d",
   173 => x"85a10481",
   174 => x"0baef40c",
   175 => x"028c050d",
   176 => x"0402fc05",
   177 => x"0d818080",
   178 => x"51c01151",
   179 => x"70fb3802",
   180 => x"84050d04",
   181 => x"02fc050d",
   182 => x"ec518371",
   183 => x"0c85c12d",
   184 => x"82710c02",
   185 => x"84050d04",
   186 => x"02f0050d",
   187 => x"805185d4",
   188 => x"2d840bec",
   189 => x"0c8be12d",
   190 => x"88a82d81",
   191 => x"f72d8352",
   192 => x"8bc62d81",
   193 => x"51848a2d",
   194 => x"ff125271",
   195 => x"8025f138",
   196 => x"840bec0c",
   197 => x"aac45185",
   198 => x"9b2da0b5",
   199 => x"2daef408",
   200 => x"802e81ef",
   201 => x"389f0bae",
   202 => x"c40c9f0b",
   203 => x"fc0cac8c",
   204 => x"518eac2d",
   205 => x"8c902d8c",
   206 => x"a32d88b4",
   207 => x"2d8ebc2d",
   208 => x"ada40b80",
   209 => x"f52dad8c",
   210 => x"0b80f52d",
   211 => x"71872b71",
   212 => x"8b2b07ad",
   213 => x"980b80f5",
   214 => x"2d708c2b",
   215 => x"7207aec4",
   216 => x"08708106",
   217 => x"53545253",
   218 => x"55555271",
   219 => x"802e8538",
   220 => x"72810753",
   221 => x"73812a70",
   222 => x"81065152",
   223 => x"71802e85",
   224 => x"38728207",
   225 => x"5373822a",
   226 => x"70810651",
   227 => x"5271802e",
   228 => x"85387284",
   229 => x"07537383",
   230 => x"2a708106",
   231 => x"51527180",
   232 => x"2e853872",
   233 => x"88075373",
   234 => x"842a7081",
   235 => x"06515271",
   236 => x"802e8538",
   237 => x"72900753",
   238 => x"73852a70",
   239 => x"81065152",
   240 => x"71802e85",
   241 => x"3872a007",
   242 => x"5373862a",
   243 => x"70810651",
   244 => x"5271802e",
   245 => x"86387280",
   246 => x"c0075373",
   247 => x"872a7081",
   248 => x"06515271",
   249 => x"802e8738",
   250 => x"7280c080",
   251 => x"07537388",
   252 => x"2a708106",
   253 => x"51527180",
   254 => x"2e873872",
   255 => x"81808007",
   256 => x"5372fc0c",
   257 => x"8652aef4",
   258 => x"08833884",
   259 => x"5271ec0c",
   260 => x"86ba0480",
   261 => x"0baef40c",
   262 => x"0290050d",
   263 => x"0471980c",
   264 => x"04ffb008",
   265 => x"aef40c04",
   266 => x"810bffb0",
   267 => x"0c04800b",
   268 => x"ffb00c04",
   269 => x"02f4050d",
   270 => x"89b604ae",
   271 => x"f40881f0",
   272 => x"2e098106",
   273 => x"8938810b",
   274 => x"aebc0c89",
   275 => x"b604aef4",
   276 => x"0881e02e",
   277 => x"09810689",
   278 => x"38810bae",
   279 => x"c00c89b6",
   280 => x"04aef408",
   281 => x"52aec008",
   282 => x"802e8838",
   283 => x"aef40881",
   284 => x"80055271",
   285 => x"842c728f",
   286 => x"065353ae",
   287 => x"bc08802e",
   288 => x"99387284",
   289 => x"29adfc05",
   290 => x"72138171",
   291 => x"2b700973",
   292 => x"0806730c",
   293 => x"51535389",
   294 => x"ac047284",
   295 => x"29adfc05",
   296 => x"72138371",
   297 => x"2b720807",
   298 => x"720c5353",
   299 => x"800baec0",
   300 => x"0c800bae",
   301 => x"bc0caf90",
   302 => x"518ab72d",
   303 => x"aef408ff",
   304 => x"24fef838",
   305 => x"800baef4",
   306 => x"0c028c05",
   307 => x"0d0402f8",
   308 => x"050dadfc",
   309 => x"528f5180",
   310 => x"72708405",
   311 => x"540cff11",
   312 => x"51708025",
   313 => x"f2380288",
   314 => x"050d0402",
   315 => x"f0050d75",
   316 => x"5188ae2d",
   317 => x"70822cfc",
   318 => x"06adfc11",
   319 => x"72109e06",
   320 => x"71087072",
   321 => x"2a708306",
   322 => x"82742b70",
   323 => x"09740676",
   324 => x"0c545156",
   325 => x"57535153",
   326 => x"88a82d71",
   327 => x"aef40c02",
   328 => x"90050d04",
   329 => x"02fc050d",
   330 => x"72518071",
   331 => x"0c800b84",
   332 => x"120c0284",
   333 => x"050d0402",
   334 => x"f0050d75",
   335 => x"70088412",
   336 => x"08535353",
   337 => x"ff547171",
   338 => x"2ea83888",
   339 => x"ae2d8413",
   340 => x"08708429",
   341 => x"14881170",
   342 => x"087081ff",
   343 => x"06841808",
   344 => x"81118706",
   345 => x"841a0c53",
   346 => x"51555151",
   347 => x"5188a82d",
   348 => x"715473ae",
   349 => x"f40c0290",
   350 => x"050d0402",
   351 => x"f4050d88",
   352 => x"ae2de008",
   353 => x"708b2a70",
   354 => x"81065152",
   355 => x"5370802e",
   356 => x"9d38af90",
   357 => x"08708429",
   358 => x"af980574",
   359 => x"81ff0671",
   360 => x"0c5151af",
   361 => x"90088111",
   362 => x"8706af90",
   363 => x"0c51728c",
   364 => x"2cbf06af",
   365 => x"b80c800b",
   366 => x"afbc0c88",
   367 => x"a12d88a8",
   368 => x"2d028c05",
   369 => x"0d0402fc",
   370 => x"050d88ae",
   371 => x"2d810baf",
   372 => x"bc0c88a8",
   373 => x"2dafbc08",
   374 => x"5170fa38",
   375 => x"0284050d",
   376 => x"0402fc05",
   377 => x"0daf9051",
   378 => x"8aa42d89",
   379 => x"ce2d8afb",
   380 => x"51889d2d",
   381 => x"0284050d",
   382 => x"0402fc05",
   383 => x"0d8fcf51",
   384 => x"85c12dff",
   385 => x"11517080",
   386 => x"25f63802",
   387 => x"84050d04",
   388 => x"02fc050d",
   389 => x"810baef0",
   390 => x"0c815184",
   391 => x"8a2d0284",
   392 => x"050d0402",
   393 => x"fc050d8c",
   394 => x"ad0488b4",
   395 => x"2d80f651",
   396 => x"89eb2dae",
   397 => x"f408f338",
   398 => x"80da5189",
   399 => x"eb2daef4",
   400 => x"08e838ae",
   401 => x"ec085189",
   402 => x"eb2daef4",
   403 => x"08dc38ae",
   404 => x"f408aef0",
   405 => x"0caef408",
   406 => x"51848a2d",
   407 => x"0284050d",
   408 => x"0402ec05",
   409 => x"0d765480",
   410 => x"52870b88",
   411 => x"1580f52d",
   412 => x"56537472",
   413 => x"248338a0",
   414 => x"53725182",
   415 => x"f82d8112",
   416 => x"8b1580f5",
   417 => x"2d545272",
   418 => x"7225de38",
   419 => x"0294050d",
   420 => x"0402f005",
   421 => x"0dafc408",
   422 => x"5481f72d",
   423 => x"800bafc8",
   424 => x"0c730880",
   425 => x"2e818038",
   426 => x"820baf88",
   427 => x"0cafc808",
   428 => x"8f06af84",
   429 => x"0c730852",
   430 => x"71832e96",
   431 => x"38718326",
   432 => x"89387181",
   433 => x"2eaf388e",
   434 => x"92047185",
   435 => x"2e9f388e",
   436 => x"92048814",
   437 => x"80f52d84",
   438 => x"1508aadc",
   439 => x"53545285",
   440 => x"9b2d7184",
   441 => x"29137008",
   442 => x"52528e96",
   443 => x"0473518c",
   444 => x"e12d8e92",
   445 => x"04aec408",
   446 => x"8815082c",
   447 => x"70810651",
   448 => x"5271802e",
   449 => x"8738aae0",
   450 => x"518e8f04",
   451 => x"aae45185",
   452 => x"9b2d8414",
   453 => x"0851859b",
   454 => x"2dafc808",
   455 => x"8105afc8",
   456 => x"0c8c1454",
   457 => x"8da10402",
   458 => x"90050d04",
   459 => x"71afc40c",
   460 => x"8d912daf",
   461 => x"c808ff05",
   462 => x"afcc0c04",
   463 => x"02e8050d",
   464 => x"afc408af",
   465 => x"d0085755",
   466 => x"80f65189",
   467 => x"eb2daef4",
   468 => x"08812a70",
   469 => x"81065152",
   470 => x"71802e9f",
   471 => x"388ee304",
   472 => x"88b42d80",
   473 => x"f65189eb",
   474 => x"2daef408",
   475 => x"f338aef0",
   476 => x"08813270",
   477 => x"aef00c51",
   478 => x"848a2d80",
   479 => x"0bafc00c",
   480 => x"8c5189eb",
   481 => x"2daef408",
   482 => x"812a7081",
   483 => x"06515271",
   484 => x"802ebd38",
   485 => x"aec808ae",
   486 => x"dc08aec8",
   487 => x"0caedc0c",
   488 => x"aecc08ae",
   489 => x"e008aecc",
   490 => x"0caee00c",
   491 => x"aed008ae",
   492 => x"e408aed0",
   493 => x"0caee40c",
   494 => x"aed408ae",
   495 => x"e808aed4",
   496 => x"0caee80c",
   497 => x"aed808ae",
   498 => x"ec08aed8",
   499 => x"0caeec0c",
   500 => x"afb808a0",
   501 => x"06528072",
   502 => x"2594388b",
   503 => x"f92d88b4",
   504 => x"2daef008",
   505 => x"813270ae",
   506 => x"f00c5184",
   507 => x"8a2daef0",
   508 => x"0881ea38",
   509 => x"aedc0851",
   510 => x"89eb2dae",
   511 => x"f408802e",
   512 => x"8938afc0",
   513 => x"088107af",
   514 => x"c00caee0",
   515 => x"085189eb",
   516 => x"2daef408",
   517 => x"802e8938",
   518 => x"afc00882",
   519 => x"07afc00c",
   520 => x"aee40851",
   521 => x"89eb2dae",
   522 => x"f408802e",
   523 => x"8938afc0",
   524 => x"088407af",
   525 => x"c00caee8",
   526 => x"085189eb",
   527 => x"2daef408",
   528 => x"802e8938",
   529 => x"afc00888",
   530 => x"07afc00c",
   531 => x"aeec0851",
   532 => x"89eb2dae",
   533 => x"f408802e",
   534 => x"8938afc0",
   535 => x"089007af",
   536 => x"c00caec8",
   537 => x"085189eb",
   538 => x"2daef408",
   539 => x"802e8a38",
   540 => x"afc00882",
   541 => x"8007afc0",
   542 => x"0caecc08",
   543 => x"5189eb2d",
   544 => x"aef40880",
   545 => x"2e8a38af",
   546 => x"c0088480",
   547 => x"07afc00c",
   548 => x"aed00851",
   549 => x"89eb2dae",
   550 => x"f408802e",
   551 => x"8a38afc0",
   552 => x"08888007",
   553 => x"afc00cae",
   554 => x"d4085189",
   555 => x"eb2daef4",
   556 => x"08802e8a",
   557 => x"38afc008",
   558 => x"908007af",
   559 => x"c00caed8",
   560 => x"085189eb",
   561 => x"2daef408",
   562 => x"802e8a38",
   563 => x"afc008a0",
   564 => x"8007afc0",
   565 => x"0cafc008",
   566 => x"ed0c98ba",
   567 => x"04aeec08",
   568 => x"5189eb2d",
   569 => x"aef40880",
   570 => x"2e8938af",
   571 => x"c0089007",
   572 => x"afc00caf",
   573 => x"c008ed0c",
   574 => x"81f55189",
   575 => x"eb2daef4",
   576 => x"08812a70",
   577 => x"81065152",
   578 => x"71a038ae",
   579 => x"dc085189",
   580 => x"eb2daef4",
   581 => x"08812a70",
   582 => x"81065152",
   583 => x"718c38af",
   584 => x"b8089006",
   585 => x"52807225",
   586 => x"bd38afb8",
   587 => x"08900652",
   588 => x"80722584",
   589 => x"388bf92d",
   590 => x"afcc0852",
   591 => x"71802e89",
   592 => x"38ff12af",
   593 => x"cc0c92e6",
   594 => x"04afc808",
   595 => x"10afc808",
   596 => x"05708429",
   597 => x"16515288",
   598 => x"1208802e",
   599 => x"8938ff51",
   600 => x"88120852",
   601 => x"712d81f2",
   602 => x"5189eb2d",
   603 => x"aef40881",
   604 => x"2a708106",
   605 => x"515271a0",
   606 => x"38aee008",
   607 => x"5189eb2d",
   608 => x"aef40881",
   609 => x"2a708106",
   610 => x"5152718c",
   611 => x"38afb808",
   612 => x"88065280",
   613 => x"7225bf38",
   614 => x"afb80888",
   615 => x"06528072",
   616 => x"2584388b",
   617 => x"f92dafc8",
   618 => x"08ff11af",
   619 => x"cc085653",
   620 => x"53737225",
   621 => x"89388114",
   622 => x"afcc0c93",
   623 => x"d6047210",
   624 => x"13708429",
   625 => x"16515288",
   626 => x"1208802e",
   627 => x"8938fe51",
   628 => x"88120852",
   629 => x"712d81fd",
   630 => x"5189eb2d",
   631 => x"aef40881",
   632 => x"2a708106",
   633 => x"51527197",
   634 => x"38aee408",
   635 => x"5189eb2d",
   636 => x"aef40881",
   637 => x"2a708106",
   638 => x"51527180",
   639 => x"2ead38af",
   640 => x"cc08802e",
   641 => x"8938800b",
   642 => x"afcc0c94",
   643 => x"ab04afc8",
   644 => x"0810afc8",
   645 => x"08057084",
   646 => x"29165152",
   647 => x"88120880",
   648 => x"2e8938fd",
   649 => x"51881208",
   650 => x"52712d81",
   651 => x"fa5189eb",
   652 => x"2daef408",
   653 => x"812a7081",
   654 => x"06515271",
   655 => x"9738aee8",
   656 => x"085189eb",
   657 => x"2daef408",
   658 => x"812a7081",
   659 => x"06515271",
   660 => x"802eae38",
   661 => x"afc808ff",
   662 => x"115452af",
   663 => x"cc087325",
   664 => x"883872af",
   665 => x"cc0c9581",
   666 => x"04711012",
   667 => x"70842916",
   668 => x"51528812",
   669 => x"08802e89",
   670 => x"38fc5188",
   671 => x"12085271",
   672 => x"2dafcc08",
   673 => x"70535473",
   674 => x"802e8a38",
   675 => x"8c15ff15",
   676 => x"55559587",
   677 => x"04820baf",
   678 => x"880c718f",
   679 => x"06af840c",
   680 => x"81eb5189",
   681 => x"eb2daef4",
   682 => x"08812a70",
   683 => x"81065152",
   684 => x"71802ead",
   685 => x"38740885",
   686 => x"2e098106",
   687 => x"a4388815",
   688 => x"80f52dff",
   689 => x"05527188",
   690 => x"1681b72d",
   691 => x"71982b52",
   692 => x"71802588",
   693 => x"38800b88",
   694 => x"1681b72d",
   695 => x"74518ce1",
   696 => x"2d81f451",
   697 => x"89eb2dae",
   698 => x"f408812a",
   699 => x"70810651",
   700 => x"5271802e",
   701 => x"b3387408",
   702 => x"852e0981",
   703 => x"06aa3888",
   704 => x"1580f52d",
   705 => x"81055271",
   706 => x"881681b7",
   707 => x"2d7181ff",
   708 => x"068b1680",
   709 => x"f52d5452",
   710 => x"72722787",
   711 => x"38728816",
   712 => x"81b72d74",
   713 => x"518ce12d",
   714 => x"80da5189",
   715 => x"eb2daef4",
   716 => x"08812a70",
   717 => x"81065152",
   718 => x"718d38af",
   719 => x"b8088106",
   720 => x"52807225",
   721 => x"81b438af",
   722 => x"c408afb8",
   723 => x"08810653",
   724 => x"53807225",
   725 => x"84388bf9",
   726 => x"2dafcc08",
   727 => x"5473802e",
   728 => x"8a388c13",
   729 => x"ff155553",
   730 => x"96dd0472",
   731 => x"08527182",
   732 => x"2ea63871",
   733 => x"82268938",
   734 => x"71812ea9",
   735 => x"3897fa04",
   736 => x"71832eb1",
   737 => x"3871842e",
   738 => x"09810680",
   739 => x"ed388813",
   740 => x"08518eac",
   741 => x"2d97fa04",
   742 => x"afcc0851",
   743 => x"88130852",
   744 => x"712d97fa",
   745 => x"04810b88",
   746 => x"14082bae",
   747 => x"c40832ae",
   748 => x"c40c97d0",
   749 => x"04881380",
   750 => x"f52d8105",
   751 => x"8b1480f5",
   752 => x"2d535471",
   753 => x"74248338",
   754 => x"80547388",
   755 => x"1481b72d",
   756 => x"8d912d97",
   757 => x"fa047508",
   758 => x"802ea238",
   759 => x"75085189",
   760 => x"eb2daef4",
   761 => x"08810652",
   762 => x"71802e8b",
   763 => x"38afcc08",
   764 => x"51841608",
   765 => x"52712d88",
   766 => x"165675da",
   767 => x"38805480",
   768 => x"0baf880c",
   769 => x"738f06af",
   770 => x"840ca052",
   771 => x"73afcc08",
   772 => x"2e098106",
   773 => x"9838afc8",
   774 => x"08ff0574",
   775 => x"32700981",
   776 => x"05707207",
   777 => x"9f2a9171",
   778 => x"31515153",
   779 => x"53715182",
   780 => x"f82d8114",
   781 => x"548e7425",
   782 => x"c638aef0",
   783 => x"08aef40c",
   784 => x"0298050d",
   785 => x"0402f405",
   786 => x"0dd45281",
   787 => x"ff720c71",
   788 => x"085381ff",
   789 => x"720c7288",
   790 => x"2b83fe80",
   791 => x"06720870",
   792 => x"81ff0651",
   793 => x"525381ff",
   794 => x"720c7271",
   795 => x"07882b72",
   796 => x"087081ff",
   797 => x"06515253",
   798 => x"81ff720c",
   799 => x"72710788",
   800 => x"2b720870",
   801 => x"81ff0672",
   802 => x"07aef40c",
   803 => x"5253028c",
   804 => x"050d0402",
   805 => x"f4050d74",
   806 => x"767181ff",
   807 => x"06d40c53",
   808 => x"53afd408",
   809 => x"85387189",
   810 => x"2b527198",
   811 => x"2ad40c71",
   812 => x"902a7081",
   813 => x"ff06d40c",
   814 => x"5171882a",
   815 => x"7081ff06",
   816 => x"d40c5171",
   817 => x"81ff06d4",
   818 => x"0c72902a",
   819 => x"7081ff06",
   820 => x"d40c51d4",
   821 => x"087081ff",
   822 => x"06515182",
   823 => x"b8bf5270",
   824 => x"81ff2e09",
   825 => x"81069438",
   826 => x"81ff0bd4",
   827 => x"0cd40870",
   828 => x"81ff06ff",
   829 => x"14545151",
   830 => x"71e53870",
   831 => x"aef40c02",
   832 => x"8c050d04",
   833 => x"02fc050d",
   834 => x"81c75181",
   835 => x"ff0bd40c",
   836 => x"ff115170",
   837 => x"8025f438",
   838 => x"0284050d",
   839 => x"0402f405",
   840 => x"0d81ff0b",
   841 => x"d40c9353",
   842 => x"805287fc",
   843 => x"80c15199",
   844 => x"932daef4",
   845 => x"088b3881",
   846 => x"ff0bd40c",
   847 => x"81539aca",
   848 => x"049a842d",
   849 => x"ff135372",
   850 => x"df3872ae",
   851 => x"f40c028c",
   852 => x"050d0402",
   853 => x"ec050d81",
   854 => x"0bafd40c",
   855 => x"8454d008",
   856 => x"708f2a70",
   857 => x"81065151",
   858 => x"5372f338",
   859 => x"72d00c9a",
   860 => x"842daae8",
   861 => x"51859b2d",
   862 => x"d008708f",
   863 => x"2a708106",
   864 => x"51515372",
   865 => x"f338810b",
   866 => x"d00cb153",
   867 => x"805284d4",
   868 => x"80c05199",
   869 => x"932daef4",
   870 => x"08812e93",
   871 => x"3872822e",
   872 => x"bd38ff13",
   873 => x"5372e538",
   874 => x"ff145473",
   875 => x"ffb0389a",
   876 => x"842d83aa",
   877 => x"52849c80",
   878 => x"c8519993",
   879 => x"2daef408",
   880 => x"812e0981",
   881 => x"06923898",
   882 => x"c52daef4",
   883 => x"0883ffff",
   884 => x"06537283",
   885 => x"aa2e9d38",
   886 => x"9a9d2d9b",
   887 => x"ef04aaf4",
   888 => x"51859b2d",
   889 => x"80539dbd",
   890 => x"04ab8c51",
   891 => x"859b2d80",
   892 => x"549d8f04",
   893 => x"81ff0bd4",
   894 => x"0cb1549a",
   895 => x"842d8fcf",
   896 => x"53805287",
   897 => x"fc80f751",
   898 => x"99932dae",
   899 => x"f40855ae",
   900 => x"f408812e",
   901 => x"0981069b",
   902 => x"3881ff0b",
   903 => x"d40c820a",
   904 => x"52849c80",
   905 => x"e9519993",
   906 => x"2daef408",
   907 => x"802e8d38",
   908 => x"9a842dff",
   909 => x"135372c9",
   910 => x"389d8204",
   911 => x"81ff0bd4",
   912 => x"0caef408",
   913 => x"5287fc80",
   914 => x"fa519993",
   915 => x"2daef408",
   916 => x"b13881ff",
   917 => x"0bd40cd4",
   918 => x"085381ff",
   919 => x"0bd40c81",
   920 => x"ff0bd40c",
   921 => x"81ff0bd4",
   922 => x"0c81ff0b",
   923 => x"d40c7286",
   924 => x"2a708106",
   925 => x"76565153",
   926 => x"729538ae",
   927 => x"f408549d",
   928 => x"8f047382",
   929 => x"2efee238",
   930 => x"ff145473",
   931 => x"feed3873",
   932 => x"afd40c73",
   933 => x"8b388152",
   934 => x"87fc80d0",
   935 => x"5199932d",
   936 => x"81ff0bd4",
   937 => x"0cd00870",
   938 => x"8f2a7081",
   939 => x"06515153",
   940 => x"72f33872",
   941 => x"d00c81ff",
   942 => x"0bd40c81",
   943 => x"5372aef4",
   944 => x"0c029405",
   945 => x"0d0402e8",
   946 => x"050d7855",
   947 => x"805681ff",
   948 => x"0bd40cd0",
   949 => x"08708f2a",
   950 => x"70810651",
   951 => x"515372f3",
   952 => x"3882810b",
   953 => x"d00c81ff",
   954 => x"0bd40c77",
   955 => x"5287fc80",
   956 => x"d1519993",
   957 => x"2d80dbc6",
   958 => x"df54aef4",
   959 => x"08802e8a",
   960 => x"38abac51",
   961 => x"859b2d9e",
   962 => x"dd0481ff",
   963 => x"0bd40cd4",
   964 => x"087081ff",
   965 => x"06515372",
   966 => x"81fe2e09",
   967 => x"81069d38",
   968 => x"80ff5398",
   969 => x"c52daef4",
   970 => x"08757084",
   971 => x"05570cff",
   972 => x"13537280",
   973 => x"25ed3881",
   974 => x"569ec204",
   975 => x"ff145473",
   976 => x"c93881ff",
   977 => x"0bd40c81",
   978 => x"ff0bd40c",
   979 => x"d008708f",
   980 => x"2a708106",
   981 => x"51515372",
   982 => x"f33872d0",
   983 => x"0c75aef4",
   984 => x"0c029805",
   985 => x"0d0402e8",
   986 => x"050d7779",
   987 => x"7b585555",
   988 => x"80537276",
   989 => x"25a33874",
   990 => x"70810556",
   991 => x"80f52d74",
   992 => x"70810556",
   993 => x"80f52d52",
   994 => x"5271712e",
   995 => x"86388151",
   996 => x"9f9b0481",
   997 => x"13539ef2",
   998 => x"04805170",
   999 => x"aef40c02",
  1000 => x"98050d04",
  1001 => x"02ec050d",
  1002 => x"76557480",
  1003 => x"2ebb389a",
  1004 => x"1580e02d",
  1005 => x"51a6a82d",
  1006 => x"aef408ae",
  1007 => x"f408b484",
  1008 => x"0caef408",
  1009 => x"5454b3e0",
  1010 => x"08802e99",
  1011 => x"38941580",
  1012 => x"e02d51a6",
  1013 => x"a82daef4",
  1014 => x"08902b83",
  1015 => x"fff00a06",
  1016 => x"70750751",
  1017 => x"5372b484",
  1018 => x"0cb48408",
  1019 => x"5372802e",
  1020 => x"9938b3d8",
  1021 => x"08fe1471",
  1022 => x"29b3ec08",
  1023 => x"05b4880c",
  1024 => x"70842bb3",
  1025 => x"e40c54a0",
  1026 => x"b004b3f0",
  1027 => x"08b4840c",
  1028 => x"b3f408b4",
  1029 => x"880cb3e0",
  1030 => x"08802e8a",
  1031 => x"38b3d808",
  1032 => x"842b53a0",
  1033 => x"ac04b3f8",
  1034 => x"08842b53",
  1035 => x"72b3e40c",
  1036 => x"0294050d",
  1037 => x"0402d805",
  1038 => x"0d800bb3",
  1039 => x"e00c8454",
  1040 => x"9ad32dae",
  1041 => x"f408802e",
  1042 => x"9538afd8",
  1043 => x"5280519d",
  1044 => x"c62daef4",
  1045 => x"08802e86",
  1046 => x"38fe54a0",
  1047 => x"e604ff14",
  1048 => x"54738024",
  1049 => x"db38738c",
  1050 => x"38abbc51",
  1051 => x"859b2d73",
  1052 => x"55a5ef04",
  1053 => x"8056810b",
  1054 => x"b48c0c88",
  1055 => x"53abd052",
  1056 => x"b08e519e",
  1057 => x"e62daef4",
  1058 => x"08762e09",
  1059 => x"81068738",
  1060 => x"aef408b4",
  1061 => x"8c0c8853",
  1062 => x"abdc52b0",
  1063 => x"aa519ee6",
  1064 => x"2daef408",
  1065 => x"8738aef4",
  1066 => x"08b48c0c",
  1067 => x"b48c0880",
  1068 => x"2e80f638",
  1069 => x"b39e0b80",
  1070 => x"f52db39f",
  1071 => x"0b80f52d",
  1072 => x"71982b71",
  1073 => x"902b07b3",
  1074 => x"a00b80f5",
  1075 => x"2d70882b",
  1076 => x"7207b3a1",
  1077 => x"0b80f52d",
  1078 => x"7107b3d6",
  1079 => x"0b80f52d",
  1080 => x"b3d70b80",
  1081 => x"f52d7188",
  1082 => x"2b07535f",
  1083 => x"54525a56",
  1084 => x"57557381",
  1085 => x"abaa2e09",
  1086 => x"81068d38",
  1087 => x"7551a5f8",
  1088 => x"2daef408",
  1089 => x"56a29504",
  1090 => x"7382d4d5",
  1091 => x"2e8738ab",
  1092 => x"e851a2d6",
  1093 => x"04afd852",
  1094 => x"75519dc6",
  1095 => x"2daef408",
  1096 => x"55aef408",
  1097 => x"802e83c7",
  1098 => x"388853ab",
  1099 => x"dc52b0aa",
  1100 => x"519ee62d",
  1101 => x"aef40889",
  1102 => x"38810bb3",
  1103 => x"e00ca2dc",
  1104 => x"048853ab",
  1105 => x"d052b08e",
  1106 => x"519ee62d",
  1107 => x"aef40880",
  1108 => x"2e8a38ab",
  1109 => x"fc51859b",
  1110 => x"2da3b604",
  1111 => x"b3d60b80",
  1112 => x"f52d5473",
  1113 => x"80d52e09",
  1114 => x"810680ca",
  1115 => x"38b3d70b",
  1116 => x"80f52d54",
  1117 => x"7381aa2e",
  1118 => x"098106ba",
  1119 => x"38800baf",
  1120 => x"d80b80f5",
  1121 => x"2d565474",
  1122 => x"81e92e83",
  1123 => x"38815474",
  1124 => x"81eb2e8c",
  1125 => x"38805573",
  1126 => x"752e0981",
  1127 => x"0682d038",
  1128 => x"afe30b80",
  1129 => x"f52d5574",
  1130 => x"8d38afe4",
  1131 => x"0b80f52d",
  1132 => x"5473822e",
  1133 => x"86388055",
  1134 => x"a5ef04af",
  1135 => x"e50b80f5",
  1136 => x"2d70b3d8",
  1137 => x"0cff05b3",
  1138 => x"dc0cafe6",
  1139 => x"0b80f52d",
  1140 => x"afe70b80",
  1141 => x"f52d5876",
  1142 => x"05778280",
  1143 => x"290570b3",
  1144 => x"e80cafe8",
  1145 => x"0b80f52d",
  1146 => x"70b3fc0c",
  1147 => x"b3e00859",
  1148 => x"57587680",
  1149 => x"2e81a338",
  1150 => x"8853abdc",
  1151 => x"52b0aa51",
  1152 => x"9ee62dae",
  1153 => x"f40881e7",
  1154 => x"38b3d808",
  1155 => x"70842bb3",
  1156 => x"e40c70b3",
  1157 => x"f80caffd",
  1158 => x"0b80f52d",
  1159 => x"affc0b80",
  1160 => x"f52d7182",
  1161 => x"802905af",
  1162 => x"fe0b80f5",
  1163 => x"2d708480",
  1164 => x"802912af",
  1165 => x"ff0b80f5",
  1166 => x"2d708180",
  1167 => x"0a291270",
  1168 => x"b4800cb3",
  1169 => x"fc087129",
  1170 => x"b3e80805",
  1171 => x"70b3ec0c",
  1172 => x"b0850b80",
  1173 => x"f52db084",
  1174 => x"0b80f52d",
  1175 => x"71828029",
  1176 => x"05b0860b",
  1177 => x"80f52d70",
  1178 => x"84808029",
  1179 => x"12b0870b",
  1180 => x"80f52d70",
  1181 => x"982b81f0",
  1182 => x"0a067205",
  1183 => x"70b3f00c",
  1184 => x"fe117e29",
  1185 => x"7705b3f4",
  1186 => x"0c525952",
  1187 => x"43545e51",
  1188 => x"5259525d",
  1189 => x"575957a5",
  1190 => x"e804afea",
  1191 => x"0b80f52d",
  1192 => x"afe90b80",
  1193 => x"f52d7182",
  1194 => x"80290570",
  1195 => x"b3e40c70",
  1196 => x"a02983ff",
  1197 => x"0570892a",
  1198 => x"70b3f80c",
  1199 => x"afef0b80",
  1200 => x"f52dafee",
  1201 => x"0b80f52d",
  1202 => x"71828029",
  1203 => x"0570b480",
  1204 => x"0c7b7129",
  1205 => x"1e70b3f4",
  1206 => x"0c7db3f0",
  1207 => x"0c7305b3",
  1208 => x"ec0c555e",
  1209 => x"51515555",
  1210 => x"80519fa4",
  1211 => x"2d815574",
  1212 => x"aef40c02",
  1213 => x"a8050d04",
  1214 => x"02f4050d",
  1215 => x"7470882a",
  1216 => x"83fe8006",
  1217 => x"7072982a",
  1218 => x"0772882b",
  1219 => x"87fc8080",
  1220 => x"0673982b",
  1221 => x"81f00a06",
  1222 => x"71730707",
  1223 => x"aef40c56",
  1224 => x"51535102",
  1225 => x"8c050d04",
  1226 => x"02f8050d",
  1227 => x"028e0580",
  1228 => x"f52d7488",
  1229 => x"2b077083",
  1230 => x"ffff06ae",
  1231 => x"f40c5102",
  1232 => x"88050d04",
  1233 => x"00ffffff",
  1234 => x"ff00ffff",
  1235 => x"ffff00ff",
  1236 => x"ffffff00",
  1237 => x"52657365",
  1238 => x"74000000",
  1239 => x"53657276",
  1240 => x"653a6175",
  1241 => x"746f6d61",
  1242 => x"7469632f",
  1243 => x"6d616e75",
  1244 => x"616c0000",
  1245 => x"42616c6c",
  1246 => x"20416e67",
  1247 => x"6c653a34",
  1248 => x"2f322061",
  1249 => x"6e676c65",
  1250 => x"73000000",
  1251 => x"42616c6c",
  1252 => x"20537065",
  1253 => x"65643a46",
  1254 => x"6173742f",
  1255 => x"536c6f77",
  1256 => x"00000000",
  1257 => x"50616464",
  1258 => x"6c652053",
  1259 => x"697a653a",
  1260 => x"736d616c",
  1261 => x"6c2f6c61",
  1262 => x"72676500",
  1263 => x"536f756e",
  1264 => x"643a4f66",
  1265 => x"662f4f6e",
  1266 => x"00000000",
  1267 => x"506c6179",
  1268 => x"6572733a",
  1269 => x"74776f2f",
  1270 => x"666f7572",
  1271 => x"00000000",
  1272 => x"4f534420",
  1273 => x"73697a65",
  1274 => x"3a73696e",
  1275 => x"676c652f",
  1276 => x"646f7562",
  1277 => x"6c650000",
  1278 => x"52616e64",
  1279 => x"6f6d2053",
  1280 => x"70656564",
  1281 => x"3a4f6666",
  1282 => x"2f4f6e00",
  1283 => x"52616e64",
  1284 => x"6f6d2041",
  1285 => x"6e676c65",
  1286 => x"3a4f6666",
  1287 => x"2f4f6e00",
  1288 => x"45786974",
  1289 => x"206d656e",
  1290 => x"75000000",
  1291 => x"4d6f6465",
  1292 => x"3a204d6f",
  1293 => x"6e6f6368",
  1294 => x"726f6d65",
  1295 => x"00000000",
  1296 => x"4d6f6465",
  1297 => x"3a204772",
  1298 => x"65797363",
  1299 => x"616c6500",
  1300 => x"4d6f6465",
  1301 => x"3a205247",
  1302 => x"42310000",
  1303 => x"4d6f6465",
  1304 => x"3a205247",
  1305 => x"42320000",
  1306 => x"4d6f6465",
  1307 => x"3a204669",
  1308 => x"656c6400",
  1309 => x"4d6f6465",
  1310 => x"3a204963",
  1311 => x"65000000",
  1312 => x"4d6f6465",
  1313 => x"3a204368",
  1314 => x"72697374",
  1315 => x"6d617300",
  1316 => x"4d6f6465",
  1317 => x"3a204d61",
  1318 => x"726b736d",
  1319 => x"616e0000",
  1320 => x"4d6f6465",
  1321 => x"3a204c61",
  1322 => x"73205665",
  1323 => x"67617300",
  1324 => x"4d6f6465",
  1325 => x"3a204159",
  1326 => x"2d332d38",
  1327 => x"35313520",
  1328 => x"636f6c6f",
  1329 => x"72730000",
  1330 => x"4d6f6465",
  1331 => x"3a205452",
  1332 => x"5120436f",
  1333 => x"6c6f7273",
  1334 => x"00000000",
  1335 => x"506c6179",
  1336 => x"65722032",
  1337 => x"3a204a6f",
  1338 => x"79737469",
  1339 => x"636b2032",
  1340 => x"00000000",
  1341 => x"506c6179",
  1342 => x"65722032",
  1343 => x"3a205061",
  1344 => x"64646c65",
  1345 => x"20656e63",
  1346 => x"6f646572",
  1347 => x"20320000",
  1348 => x"506c6179",
  1349 => x"65722031",
  1350 => x"3a204a6f",
  1351 => x"79737469",
  1352 => x"636b2031",
  1353 => x"00000000",
  1354 => x"506c6179",
  1355 => x"65722031",
  1356 => x"3a205061",
  1357 => x"64646c65",
  1358 => x"20656e63",
  1359 => x"6f646572",
  1360 => x"20310000",
  1361 => x"496e6974",
  1362 => x"69616c69",
  1363 => x"7a696e67",
  1364 => x"20534420",
  1365 => x"63617264",
  1366 => x"0a000000",
  1367 => x"16200000",
  1368 => x"14200000",
  1369 => x"15200000",
  1370 => x"53442069",
  1371 => x"6e69742e",
  1372 => x"2e2e0a00",
  1373 => x"53442063",
  1374 => x"61726420",
  1375 => x"72657365",
  1376 => x"74206661",
  1377 => x"696c6564",
  1378 => x"210a0000",
  1379 => x"53444843",
  1380 => x"20657272",
  1381 => x"6f72210a",
  1382 => x"00000000",
  1383 => x"57726974",
  1384 => x"65206661",
  1385 => x"696c6564",
  1386 => x"0a000000",
  1387 => x"52656164",
  1388 => x"20666169",
  1389 => x"6c65640a",
  1390 => x"00000000",
  1391 => x"43617264",
  1392 => x"20696e69",
  1393 => x"74206661",
  1394 => x"696c6564",
  1395 => x"0a000000",
  1396 => x"46415431",
  1397 => x"36202020",
  1398 => x"00000000",
  1399 => x"46415433",
  1400 => x"32202020",
  1401 => x"00000000",
  1402 => x"4e6f2070",
  1403 => x"61727469",
  1404 => x"74696f6e",
  1405 => x"20736967",
  1406 => x"0a000000",
  1407 => x"42616420",
  1408 => x"70617274",
  1409 => x"0a000000",
  1410 => x"00000002",
  1411 => x"00000002",
  1412 => x"00001354",
  1413 => x"000002d4",
  1414 => x"00000001",
  1415 => x"0000135c",
  1416 => x"00000000",
  1417 => x"00000001",
  1418 => x"00001374",
  1419 => x"00000001",
  1420 => x"00000001",
  1421 => x"0000138c",
  1422 => x"00000002",
  1423 => x"00000001",
  1424 => x"000013a4",
  1425 => x"00000003",
  1426 => x"00000001",
  1427 => x"000013bc",
  1428 => x"00000004",
  1429 => x"00000001",
  1430 => x"000013cc",
  1431 => x"00000006",
  1432 => x"00000001",
  1433 => x"000013e0",
  1434 => x"00000005",
  1435 => x"00000001",
  1436 => x"000013f8",
  1437 => x"00000007",
  1438 => x"00000001",
  1439 => x"0000140c",
  1440 => x"00000008",
  1441 => x"00000003",
  1442 => x"000016f4",
  1443 => x"00000002",
  1444 => x"00000003",
  1445 => x"000016ec",
  1446 => x"00000002",
  1447 => x"00000003",
  1448 => x"000016c0",
  1449 => x"0000000b",
  1450 => x"00000002",
  1451 => x"00001420",
  1452 => x"00000623",
  1453 => x"00000000",
  1454 => x"00000000",
  1455 => x"00000000",
  1456 => x"0000142c",
  1457 => x"00001440",
  1458 => x"00001450",
  1459 => x"0000145c",
  1460 => x"00001468",
  1461 => x"00001474",
  1462 => x"00001480",
  1463 => x"00001490",
  1464 => x"000014a0",
  1465 => x"000014b0",
  1466 => x"000014c8",
  1467 => x"000014dc",
  1468 => x"000014f4",
  1469 => x"00001510",
  1470 => x"00001528",
  1471 => x"00000000",
  1472 => x"00000000",
  1473 => x"00000000",
  1474 => x"00000000",
  1475 => x"00000000",
  1476 => x"00000000",
  1477 => x"00000000",
  1478 => x"00000000",
  1479 => x"00000000",
  1480 => x"00000000",
  1481 => x"00000000",
  1482 => x"00000000",
  1483 => x"00000000",
  1484 => x"00000000",
  1485 => x"00000000",
  1486 => x"00000000",
  1487 => x"00000000",
  1488 => x"00000000",
  1489 => x"00000006",
  1490 => x"00000043",
  1491 => x"00000042",
  1492 => x"0000003b",
  1493 => x"0000004b",
  1494 => x"0000007e",
  1495 => x"00000003",
  1496 => x"0000000b",
  1497 => x"00000083",
  1498 => x"00000023",
  1499 => x"0000007e",
  1500 => x"00000000",
	others => x"00000000"
);

begin

process (clk)
begin
	if (clk'event and clk = '1') then
		if (from_zpu.memAWriteEnable = '1') and (from_zpu.memBWriteEnable = '1') and (from_zpu.memAAddr=from_zpu.memBAddr) and (from_zpu.memAWrite/=from_zpu.memBWrite) then
			report "write collision" severity failure;
		end if;
	
		if (from_zpu.memAWriteEnable = '1') then
			ram(to_integer(unsigned(from_zpu.memAAddr(maxAddrBitBRAM downto 2)))) := from_zpu.memAWrite;
			to_zpu.memARead <= from_zpu.memAWrite;
		else
			to_zpu.memARead <= ram(to_integer(unsigned(from_zpu.memAAddr(maxAddrBitBRAM downto 2))));
		end if;
	end if;
end process;

process (clk)
begin
	if (clk'event and clk = '1') then
		if (from_zpu.memBWriteEnable = '1') then
			ram(to_integer(unsigned(from_zpu.memBAddr(maxAddrBitBRAM downto 2)))) := from_zpu.memBWrite;
			to_zpu.memBRead <= from_zpu.memBWrite;
		else
			to_zpu.memBRead <= ram(to_integer(unsigned(from_zpu.memBAddr(maxAddrBitBRAM downto 2))));
		end if;
	end if;
end process;


end arch;

