12
1e
31
2e
30
30
20
4b
2e
76
2e
53
65
6e
67
62
75
73
63
68
20
32
34
2f
34
2d
27
39
34
00
00
ff
65
32
66
32
67
28
83
50
84
60
62
64
69
00
6a
01
6b
00
00
c1
22
b0
60
01
82
05
60
28
52
00
12
32
a3
38
d3
48
a3
38
d3
48
00
c1
d5
68
3f
00
12
78
22
b0
60
01
32
00
82
05
22
ec
83
50
84
60
60
07
e0
a1
22
94
60
08
e0
a1
22
8c
c0
03
40
00
22
9e
c0
03
40
00
22
a6
12
44
80
b0
70
03
80
06
80
06
f0
30
80
70
70
11
61
1b
d0
1a
12
8a
75
01
45
6e
65
6d
00
ee
60
01
85
05
4f
00
65
00
00
ee
77
01
47
46
67
45
00
ee
60
01
87
05
47
14
67
15
00
ee
80
90
61
2d
81
05
88
10
61
00
80
70
a3
2c
d0
11
80
84
61
00
d0
11
7a
01
4a
04
6a
01
4a
01
a3
2e
4a
02
a3
30
4a
03
a3
32
61
00
60
00
d0
11
60
08
d0
11
60
70
d0
11
60
78
d0
11
00
ee
32
00
00
ee
c0
0f
80
74
70
08
61
00
a3
38
62
2d
4b
1e
23
10
3b
21
d0
18
7b
01
80
90
82
05
39
0b
79
01
00
ee
7b
03
a3
34
80
70
70
05
d0
11
70
08
d0
11
70
08
d0
11
70
08
a3
36
d0
11
62
64
00
ee
88
00
88
00
55
00
22
00
ff
00
f8
00
db
ff
db
18
24
e7
e7
db
