-- ZPU
--
-- Copyright 2004-2008 oharboe - �yvind Harboe - oyvind.harboe@zylin.com
-- Modified by Alastair M. Robinson for the ZPUFlex project.
--
-- The FreeBSD license
-- 
-- Redistribution and use in source and binary forms, with or without
-- modification, are permitted provided that the following conditions
-- are met:
-- 
-- 1. Redistributions of source code must retain the above copyright
--    notice, this list of conditions and the following disclaimer.
-- 2. Redistributions in binary form must reproduce the above
--    copyright notice, this list of conditions and the following
--    disclaimer in the documentation and/or other materials
--    provided with the distribution.
-- 
-- THIS SOFTWARE IS PROVIDED BY THE ZPU PROJECT ``AS IS'' AND ANY
-- EXPRESS OR IMPLIED WARRANTIES, INCLUDING, BUT NOT LIMITED TO,
-- THE IMPLIED WARRANTIES OF MERCHANTABILITY AND FITNESS FOR A
-- PARTICULAR PURPOSE ARE DISCLAIMED. IN NO EVENT SHALL THE
-- ZPU PROJECT OR CONTRIBUTORS BE LIABLE FOR ANY DIRECT,
-- INDIRECT, INCIDENTAL, SPECIAL, EXEMPLARY, OR CONSEQUENTIAL DAMAGES
-- (INCLUDING, BUT NOT LIMITED TO, PROCUREMENT OF SUBSTITUTE GOODS
-- OR SERVICES; LOSS OF USE, DATA, OR PROFITS; OR BUSINESS INTERRUPTION)
-- HOWEVER CAUSED AND ON ANY THEORY OF LIABILITY, WHETHER IN CONTRACT,
-- STRICT LIABILITY, OR TORT (INCLUDING NEGLIGENCE OR OTHERWISE)
-- ARISING IN ANY WAY OUT OF THE USE OF THIS SOFTWARE, EVEN IF
-- ADVISED OF THE POSSIBILITY OF SUCH DAMAGE.
-- 
-- The views and conclusions contained in the software and documentation
-- are those of the authors and should not be interpreted as representing
-- official policies, either expressed or implied, of the ZPU Project.

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;


library work;
use work.zpupkg.all;

entity CtrlROM_ROM is
generic
	(
		maxAddrBitBRAM : integer := maxAddrBitBRAMLimit -- Specify your actual ROM size to save LEs and unnecessary block RAM usage.
	);
port (
	clk : in std_logic;
	areset : in std_logic := '0';
	from_zpu : in ZPU_ToROM;
	to_zpu : out ZPU_FromROM
);
end CtrlROM_ROM;

architecture arch of CtrlROM_ROM is

type ram_type is array(natural range 0 to ((2**(maxAddrBitBRAM+1))/4)-1) of std_logic_vector(wordSize-1 downto 0);

shared variable ram : ram_type :=
(
     0 => x"0b0b0b0b",
     1 => x"8c0b0b0b",
     2 => x"0b81e004",
     3 => x"0b0b0b0b",
     4 => x"8c04ff0d",
     5 => x"80040400",
     6 => x"00000016",
     7 => x"00000000",
     8 => x"0b0b80cb",
     9 => x"f4080b0b",
    10 => x"80cbf808",
    11 => x"0b0b80cb",
    12 => x"fc080b0b",
    13 => x"0b0b9808",
    14 => x"2d0b0b80",
    15 => x"cbfc0c0b",
    16 => x"0b80cbf8",
    17 => x"0c0b0b80",
    18 => x"cbf40c04",
    19 => x"00000000",
    20 => x"00000000",
    21 => x"00000000",
    22 => x"00000000",
    23 => x"00000000",
    24 => x"71fd0608",
    25 => x"72830609",
    26 => x"81058205",
    27 => x"832b2a83",
    28 => x"ffff0652",
    29 => x"0471fc06",
    30 => x"08728306",
    31 => x"09810583",
    32 => x"05101010",
    33 => x"2a81ff06",
    34 => x"520471fd",
    35 => x"060883ff",
    36 => x"ff738306",
    37 => x"09810582",
    38 => x"05832b2b",
    39 => x"09067383",
    40 => x"ffff0673",
    41 => x"83060981",
    42 => x"05820583",
    43 => x"2b0b2b07",
    44 => x"72fc060c",
    45 => x"51510471",
    46 => x"fc06080b",
    47 => x"0b80c3d4",
    48 => x"73830610",
    49 => x"10050806",
    50 => x"7381ff06",
    51 => x"73830609",
    52 => x"81058305",
    53 => x"1010102b",
    54 => x"0772fc06",
    55 => x"0c515104",
    56 => x"80cbf470",
    57 => x"80d6a827",
    58 => x"8b388071",
    59 => x"70840553",
    60 => x"0c81e304",
    61 => x"8c519691",
    62 => x"0402fc05",
    63 => x"0df88051",
    64 => x"8f0b80cc",
    65 => x"840c9f0b",
    66 => x"80cc880c",
    67 => x"a0717081",
    68 => x"05533480",
    69 => x"cc8808ff",
    70 => x"0580cc88",
    71 => x"0c80cc88",
    72 => x"088025e8",
    73 => x"3880cc84",
    74 => x"08ff0580",
    75 => x"cc840c80",
    76 => x"cc840880",
    77 => x"25d03880",
    78 => x"0b80cc88",
    79 => x"0c800b80",
    80 => x"cc840c02",
    81 => x"84050d04",
    82 => x"02f0050d",
    83 => x"f88053f8",
    84 => x"a05483bf",
    85 => x"52737081",
    86 => x"05553351",
    87 => x"70737081",
    88 => x"055534ff",
    89 => x"12527180",
    90 => x"25eb38fb",
    91 => x"c0539f52",
    92 => x"a0737081",
    93 => x"055534ff",
    94 => x"12527180",
    95 => x"25f23802",
    96 => x"90050d04",
    97 => x"02f4050d",
    98 => x"74538e0b",
    99 => x"80cc8408",
   100 => x"25913882",
   101 => x"c82d80cc",
   102 => x"8408ff05",
   103 => x"80cc840c",
   104 => x"838a0480",
   105 => x"cc840880",
   106 => x"cc880853",
   107 => x"51728a2e",
   108 => x"098106be",
   109 => x"38715171",
   110 => x"9f24a438",
   111 => x"80cc8408",
   112 => x"a02911f8",
   113 => x"80115151",
   114 => x"a0713480",
   115 => x"cc880881",
   116 => x"0580cc88",
   117 => x"0c80cc88",
   118 => x"08519f71",
   119 => x"25de3880",
   120 => x"0b80cc88",
   121 => x"0c80cc84",
   122 => x"08810580",
   123 => x"cc840c84",
   124 => x"880470a0",
   125 => x"2912f880",
   126 => x"11515172",
   127 => x"713480cc",
   128 => x"88088105",
   129 => x"80cc880c",
   130 => x"80cc8808",
   131 => x"a02e0981",
   132 => x"06913880",
   133 => x"0b80cc88",
   134 => x"0c80cc84",
   135 => x"08810580",
   136 => x"cc840c02",
   137 => x"8c050d04",
   138 => x"02e8050d",
   139 => x"77795656",
   140 => x"880bfc16",
   141 => x"77712c8f",
   142 => x"06545254",
   143 => x"80537272",
   144 => x"25953871",
   145 => x"53fbe014",
   146 => x"51877134",
   147 => x"8114ff14",
   148 => x"545472f1",
   149 => x"387153f9",
   150 => x"1576712c",
   151 => x"87065351",
   152 => x"71802e8b",
   153 => x"38fbe014",
   154 => x"51717134",
   155 => x"81145472",
   156 => x"8e249538",
   157 => x"8f733153",
   158 => x"fbe01451",
   159 => x"a0713481",
   160 => x"14ff1454",
   161 => x"5472f138",
   162 => x"0298050d",
   163 => x"0402ec05",
   164 => x"0d800b80",
   165 => x"cc8c0cf6",
   166 => x"8c08f690",
   167 => x"0871882c",
   168 => x"565481ff",
   169 => x"06527372",
   170 => x"25893871",
   171 => x"54820b80",
   172 => x"cc8c0c72",
   173 => x"882c7381",
   174 => x"ff065455",
   175 => x"7473258d",
   176 => x"387280cc",
   177 => x"8c088407",
   178 => x"80cc8c0c",
   179 => x"5573842b",
   180 => x"86a07125",
   181 => x"83713170",
   182 => x"0b0b80c7",
   183 => x"d80c8171",
   184 => x"2bff05f6",
   185 => x"880cfc08",
   186 => x"fea414ff",
   187 => x"132c7988",
   188 => x"29fed005",
   189 => x"70812c80",
   190 => x"cc8c0852",
   191 => x"59535155",
   192 => x"51525476",
   193 => x"802e8538",
   194 => x"70810751",
   195 => x"70f6940c",
   196 => x"71098105",
   197 => x"f6800c72",
   198 => x"098105f6",
   199 => x"840c0294",
   200 => x"050d0402",
   201 => x"f4050d74",
   202 => x"53727081",
   203 => x"055480f5",
   204 => x"2d527180",
   205 => x"2e893871",
   206 => x"5183842d",
   207 => x"86a90481",
   208 => x"0b80cbf4",
   209 => x"0c028c05",
   210 => x"0d0402fc",
   211 => x"050d8180",
   212 => x"8051c011",
   213 => x"5170fb38",
   214 => x"0284050d",
   215 => x"0402fc05",
   216 => x"0dec5183",
   217 => x"710c86ca",
   218 => x"2d82710c",
   219 => x"0284050d",
   220 => x"0486ca2d",
   221 => x"86ca2d86",
   222 => x"ca2d86ca",
   223 => x"2d86ca2d",
   224 => x"86ca2d86",
   225 => x"ca2d86ca",
   226 => x"2d86ca2d",
   227 => x"86ca2d86",
   228 => x"ca2d86ca",
   229 => x"2d86ca2d",
   230 => x"86ca2d86",
   231 => x"ca2d86ca",
   232 => x"2d86ca2d",
   233 => x"86ca2d86",
   234 => x"ca2d86ca",
   235 => x"2d86ca2d",
   236 => x"86ca2d86",
   237 => x"ca2d86ca",
   238 => x"2d86ca2d",
   239 => x"86ca2d86",
   240 => x"ca2d86ca",
   241 => x"2d86ca2d",
   242 => x"86ca2d86",
   243 => x"ca2d86ca",
   244 => x"2d86ca2d",
   245 => x"86ca2d86",
   246 => x"ca2d86ca",
   247 => x"2d86ca2d",
   248 => x"86ca2d86",
   249 => x"ca2d86ca",
   250 => x"2d86ca2d",
   251 => x"86ca2d86",
   252 => x"ca2d86ca",
   253 => x"2d86ca2d",
   254 => x"86ca2d86",
   255 => x"ca2d86ca",
   256 => x"2d86ca2d",
   257 => x"86ca2d86",
   258 => x"ca2d86ca",
   259 => x"2d86ca2d",
   260 => x"86ca2d86",
   261 => x"ca2d86ca",
   262 => x"2d86ca2d",
   263 => x"86ca2d86",
   264 => x"ca2d86ca",
   265 => x"2d86ca2d",
   266 => x"86ca2d86",
   267 => x"ca2d86ca",
   268 => x"2d86ca2d",
   269 => x"86ca2d86",
   270 => x"ca2d86ca",
   271 => x"2d86ca2d",
   272 => x"86ca2d86",
   273 => x"ca2d86ca",
   274 => x"2d86ca2d",
   275 => x"86ca2d86",
   276 => x"ca2d86ca",
   277 => x"2d86ca2d",
   278 => x"86ca2d86",
   279 => x"ca2d86ca",
   280 => x"2d86ca2d",
   281 => x"86ca2d86",
   282 => x"ca2d86ca",
   283 => x"2d86ca2d",
   284 => x"86ca2d86",
   285 => x"ca2d86ca",
   286 => x"2d86ca2d",
   287 => x"86ca2d86",
   288 => x"ca2d86ca",
   289 => x"2d86ca2d",
   290 => x"86ca2d86",
   291 => x"ca2d86ca",
   292 => x"2d86ca2d",
   293 => x"86ca2d86",
   294 => x"ca2d86ca",
   295 => x"2d86ca2d",
   296 => x"86ca2d86",
   297 => x"ca2d86ca",
   298 => x"2d86ca2d",
   299 => x"86ca2d86",
   300 => x"ca2d86ca",
   301 => x"2d86ca2d",
   302 => x"86ca2d86",
   303 => x"ca2d86ca",
   304 => x"2d86ca2d",
   305 => x"86ca2d86",
   306 => x"ca2d86ca",
   307 => x"2d86ca2d",
   308 => x"86ca2d86",
   309 => x"ca2d86ca",
   310 => x"2d86ca2d",
   311 => x"86ca2d86",
   312 => x"ca2d86ca",
   313 => x"2d86ca2d",
   314 => x"86ca2d86",
   315 => x"ca2d86ca",
   316 => x"2d86ca2d",
   317 => x"86ca2d86",
   318 => x"ca2d86ca",
   319 => x"2d86ca2d",
   320 => x"86ca2d86",
   321 => x"ca2d86ca",
   322 => x"2d86ca2d",
   323 => x"86ca2d86",
   324 => x"ca2d86ca",
   325 => x"2d86ca2d",
   326 => x"86ca2d86",
   327 => x"ca2d86ca",
   328 => x"2d86ca2d",
   329 => x"86ca2d86",
   330 => x"ca2d86ca",
   331 => x"2d86ca2d",
   332 => x"86ca2d86",
   333 => x"ca2d86ca",
   334 => x"2d86ca2d",
   335 => x"86ca2d86",
   336 => x"ca2d86ca",
   337 => x"2d86ca2d",
   338 => x"86ca2d86",
   339 => x"ca2d86ca",
   340 => x"2d86ca2d",
   341 => x"86ca2d86",
   342 => x"ca2d86ca",
   343 => x"2d86ca2d",
   344 => x"86ca2d86",
   345 => x"ca2d86ca",
   346 => x"2d86ca2d",
   347 => x"86ca2d86",
   348 => x"ca2d86ca",
   349 => x"2d86ca2d",
   350 => x"86ca2d86",
   351 => x"ca2d86ca",
   352 => x"2d86ca2d",
   353 => x"86ca2d86",
   354 => x"ca2d86ca",
   355 => x"2d86ca2d",
   356 => x"86ca2d86",
   357 => x"ca2d86ca",
   358 => x"2d86ca2d",
   359 => x"86ca2d86",
   360 => x"ca2d86ca",
   361 => x"2d86ca2d",
   362 => x"86ca2d86",
   363 => x"ca2d86ca",
   364 => x"2d86ca2d",
   365 => x"86ca2d86",
   366 => x"ca2d86ca",
   367 => x"2d86ca2d",
   368 => x"86ca2d86",
   369 => x"ca2d86ca",
   370 => x"2d86ca2d",
   371 => x"86ca2d86",
   372 => x"ca2d86ca",
   373 => x"2d86ca2d",
   374 => x"86ca2d86",
   375 => x"ca2d86ca",
   376 => x"2d86ca2d",
   377 => x"86ca2d86",
   378 => x"ca2d86ca",
   379 => x"2d86ca2d",
   380 => x"86ca2d86",
   381 => x"ca2d86ca",
   382 => x"2d86ca2d",
   383 => x"86ca2d86",
   384 => x"ca2d86ca",
   385 => x"2d86ca2d",
   386 => x"86ca2d86",
   387 => x"ca2d86ca",
   388 => x"2d86ca2d",
   389 => x"86ca2d86",
   390 => x"ca2d86ca",
   391 => x"2d86ca2d",
   392 => x"86ca2d86",
   393 => x"ca2d86ca",
   394 => x"2d86ca2d",
   395 => x"86ca2d86",
   396 => x"ca2d86ca",
   397 => x"2d86ca2d",
   398 => x"86ca2d86",
   399 => x"ca2d86ca",
   400 => x"2d86ca2d",
   401 => x"86ca2d86",
   402 => x"ca2d86ca",
   403 => x"2d86ca2d",
   404 => x"86ca2d86",
   405 => x"ca2d86ca",
   406 => x"2d86ca2d",
   407 => x"86ca2d86",
   408 => x"ca2d86ca",
   409 => x"2d86ca2d",
   410 => x"86ca2d86",
   411 => x"ca2d86ca",
   412 => x"2d86ca2d",
   413 => x"86ca2d86",
   414 => x"ca2d86ca",
   415 => x"2d86ca2d",
   416 => x"86ca2d86",
   417 => x"ca2d86ca",
   418 => x"2d86ca2d",
   419 => x"86ca2d86",
   420 => x"ca2d86ca",
   421 => x"2d86ca2d",
   422 => x"86ca2d86",
   423 => x"ca2d86ca",
   424 => x"2d86ca2d",
   425 => x"86ca2d86",
   426 => x"ca2d86ca",
   427 => x"2d86ca2d",
   428 => x"86ca2d86",
   429 => x"ca2d86ca",
   430 => x"2d86ca2d",
   431 => x"86ca2d86",
   432 => x"ca2d86ca",
   433 => x"2d86ca2d",
   434 => x"86ca2d86",
   435 => x"ca2d86ca",
   436 => x"2d86ca2d",
   437 => x"86ca2d86",
   438 => x"ca2d86ca",
   439 => x"2d86ca2d",
   440 => x"86ca2d86",
   441 => x"ca2d86ca",
   442 => x"2d86ca2d",
   443 => x"86ca2d86",
   444 => x"ca2d86ca",
   445 => x"2d86ca2d",
   446 => x"86ca2d86",
   447 => x"ca2d86ca",
   448 => x"2d86ca2d",
   449 => x"86ca2d86",
   450 => x"ca2d86ca",
   451 => x"2d86ca2d",
   452 => x"86ca2d86",
   453 => x"ca2d86ca",
   454 => x"2d86ca2d",
   455 => x"86ca2d86",
   456 => x"ca2d86ca",
   457 => x"2d86ca2d",
   458 => x"86ca2d86",
   459 => x"ca2d86ca",
   460 => x"2d86ca2d",
   461 => x"86ca2d86",
   462 => x"ca2d86ca",
   463 => x"2d86ca2d",
   464 => x"86ca2d86",
   465 => x"ca2d86ca",
   466 => x"2d86ca2d",
   467 => x"86ca2d86",
   468 => x"ca2d86ca",
   469 => x"2d86ca2d",
   470 => x"86ca2d86",
   471 => x"ca2d86ca",
   472 => x"2d86ca2d",
   473 => x"86ca2d86",
   474 => x"ca2d86ca",
   475 => x"2d86ca2d",
   476 => x"86ca2d86",
   477 => x"ca2d86ca",
   478 => x"2d86ca2d",
   479 => x"86ca2d86",
   480 => x"ca2d86ca",
   481 => x"2d86ca2d",
   482 => x"86ca2d86",
   483 => x"ca2d86ca",
   484 => x"2d86ca2d",
   485 => x"86ca2d86",
   486 => x"ca2d86ca",
   487 => x"2d86ca2d",
   488 => x"86ca2d86",
   489 => x"ca2d86ca",
   490 => x"2d86ca2d",
   491 => x"86ca2d86",
   492 => x"ca2d86ca",
   493 => x"2d86ca2d",
   494 => x"86ca2d86",
   495 => x"ca2d86ca",
   496 => x"2d86ca2d",
   497 => x"86ca2d86",
   498 => x"ca2d86ca",
   499 => x"2d86ca2d",
   500 => x"86ca2d86",
   501 => x"ca2d86ca",
   502 => x"2d86ca2d",
   503 => x"86ca2d86",
   504 => x"ca2d86ca",
   505 => x"2d86ca2d",
   506 => x"86ca2d86",
   507 => x"ca2d86ca",
   508 => x"2d86ca2d",
   509 => x"86ca2d86",
   510 => x"ca2d86ca",
   511 => x"2d86ca2d",
   512 => x"86ca2d86",
   513 => x"ca2d86ca",
   514 => x"2d86ca2d",
   515 => x"86ca2d86",
   516 => x"ca2d86ca",
   517 => x"2d86ca2d",
   518 => x"86ca2d86",
   519 => x"ca2d86ca",
   520 => x"2d86ca2d",
   521 => x"86ca2d86",
   522 => x"ca2d86ca",
   523 => x"2d86ca2d",
   524 => x"86ca2d86",
   525 => x"ca2d86ca",
   526 => x"2d86ca2d",
   527 => x"86ca2d86",
   528 => x"ca2d86ca",
   529 => x"2d86ca2d",
   530 => x"86ca2d86",
   531 => x"ca2d86ca",
   532 => x"2d86ca2d",
   533 => x"86ca2d86",
   534 => x"ca2d86ca",
   535 => x"2d86ca2d",
   536 => x"86ca2d86",
   537 => x"ca2d86ca",
   538 => x"2d86ca2d",
   539 => x"86ca2d86",
   540 => x"ca2d86ca",
   541 => x"2d86ca2d",
   542 => x"86ca2d86",
   543 => x"ca2d86ca",
   544 => x"2d86ca2d",
   545 => x"86ca2d86",
   546 => x"ca2d86ca",
   547 => x"2d86ca2d",
   548 => x"86ca2d86",
   549 => x"ca2d86ca",
   550 => x"2d86ca2d",
   551 => x"86ca2d86",
   552 => x"ca2d86ca",
   553 => x"2d86ca2d",
   554 => x"86ca2d86",
   555 => x"ca2d86ca",
   556 => x"2d86ca2d",
   557 => x"86ca2d86",
   558 => x"ca2d86ca",
   559 => x"2d86ca2d",
   560 => x"86ca2d86",
   561 => x"ca2d86ca",
   562 => x"2d86ca2d",
   563 => x"86ca2d86",
   564 => x"ca2d86ca",
   565 => x"2d86ca2d",
   566 => x"86ca2d86",
   567 => x"ca2d86ca",
   568 => x"2d86ca2d",
   569 => x"86ca2d86",
   570 => x"ca2d86ca",
   571 => x"2d86ca2d",
   572 => x"86ca2d86",
   573 => x"ca2d86ca",
   574 => x"2d86ca2d",
   575 => x"86ca2d86",
   576 => x"ca2d86ca",
   577 => x"2d86ca2d",
   578 => x"86ca2d86",
   579 => x"ca2d86ca",
   580 => x"2d86ca2d",
   581 => x"86ca2d86",
   582 => x"ca2d86ca",
   583 => x"2d86ca2d",
   584 => x"86ca2d86",
   585 => x"ca2d86ca",
   586 => x"2d86ca2d",
   587 => x"86ca2d86",
   588 => x"ca2d86ca",
   589 => x"2d86ca2d",
   590 => x"86ca2d86",
   591 => x"ca2d86ca",
   592 => x"2d86ca2d",
   593 => x"86ca2d86",
   594 => x"ca2d86ca",
   595 => x"2d86ca2d",
   596 => x"86ca2d86",
   597 => x"ca2d86ca",
   598 => x"2d86ca2d",
   599 => x"86ca2d86",
   600 => x"ca2d86ca",
   601 => x"2d86ca2d",
   602 => x"86ca2d86",
   603 => x"ca2d86ca",
   604 => x"2d86ca2d",
   605 => x"86ca2d86",
   606 => x"ca2d86ca",
   607 => x"2d86ca2d",
   608 => x"86ca2d86",
   609 => x"ca2d86ca",
   610 => x"2d86ca2d",
   611 => x"86ca2d86",
   612 => x"ca2d86ca",
   613 => x"2d86ca2d",
   614 => x"86ca2d86",
   615 => x"ca2d86ca",
   616 => x"2d86ca2d",
   617 => x"86ca2d86",
   618 => x"ca2d86ca",
   619 => x"2d86ca2d",
   620 => x"86ca2d86",
   621 => x"ca2d86ca",
   622 => x"2d86ca2d",
   623 => x"86ca2d86",
   624 => x"ca2d86ca",
   625 => x"2d86ca2d",
   626 => x"86ca2d86",
   627 => x"ca2d86ca",
   628 => x"2d86ca2d",
   629 => x"86ca2d86",
   630 => x"ca2d86ca",
   631 => x"2d86ca2d",
   632 => x"86ca2d86",
   633 => x"ca2d86ca",
   634 => x"2d86ca2d",
   635 => x"86ca2d86",
   636 => x"ca2d86ca",
   637 => x"2d86ca2d",
   638 => x"86ca2d86",
   639 => x"ca2d86ca",
   640 => x"2d86ca2d",
   641 => x"86ca2d86",
   642 => x"ca2d86ca",
   643 => x"2d86ca2d",
   644 => x"86ca2d86",
   645 => x"ca2d86ca",
   646 => x"2d86ca2d",
   647 => x"86ca2d86",
   648 => x"ca2d86ca",
   649 => x"2d86ca2d",
   650 => x"86ca2d86",
   651 => x"ca2d86ca",
   652 => x"2d0402dc",
   653 => x"050d7a53",
   654 => x"8059840b",
   655 => x"ec0c7252",
   656 => x"80cc9051",
   657 => x"bab62d80",
   658 => x"cbf40879",
   659 => x"2e819d38",
   660 => x"80cc9408",
   661 => x"79ff1256",
   662 => x"59557485",
   663 => x"2e098106",
   664 => x"a4387251",
   665 => x"86a32d86",
   666 => x"f12d86f1",
   667 => x"2d86f12d",
   668 => x"86f12d86",
   669 => x"f12d86f1",
   670 => x"2d80c7dc",
   671 => x"519ea42d",
   672 => x"81539687",
   673 => x"0473802e",
   674 => x"8b388118",
   675 => x"74812a55",
   676 => x"58958504",
   677 => x"f7185881",
   678 => x"59807525",
   679 => x"80ce3877",
   680 => x"52735184",
   681 => x"a82d80cc",
   682 => x"e05280cc",
   683 => x"9051bd83",
   684 => x"2d80cbf4",
   685 => x"08802e9b",
   686 => x"3880cce0",
   687 => x"5783fc56",
   688 => x"76708405",
   689 => x"5808e80c",
   690 => x"fc165675",
   691 => x"8025f138",
   692 => x"95db0480",
   693 => x"cbf40859",
   694 => x"84805580",
   695 => x"cc9051bc",
   696 => x"d32dfc80",
   697 => x"15811555",
   698 => x"55959904",
   699 => x"80cc9408",
   700 => x"f80c7880",
   701 => x"2e883880",
   702 => x"c8bc5196",
   703 => x"820480c8",
   704 => x"98519ea4",
   705 => x"2d785372",
   706 => x"80cbf40c",
   707 => x"02a4050d",
   708 => x"0402f005",
   709 => x"0d805186",
   710 => x"dd2d840b",
   711 => x"ec0c9bd3",
   712 => x"2d98882d",
   713 => x"81f92d83",
   714 => x"529bb62d",
   715 => x"8151858d",
   716 => x"2dff1252",
   717 => x"718025f1",
   718 => x"38840bec",
   719 => x"0c80c68c",
   720 => x"5186a32d",
   721 => x"b0ee2d80",
   722 => x"cbf40880",
   723 => x"2e81a238",
   724 => x"810bec0c",
   725 => x"840bec0c",
   726 => x"94b25180",
   727 => x"c3cc2d80",
   728 => x"c7dc519e",
   729 => x"a42d9bf5",
   730 => x"2d98942d",
   731 => x"9eb72d80",
   732 => x"c7f00b80",
   733 => x"f52d80ca",
   734 => x"88087081",
   735 => x"06545553",
   736 => x"71802e85",
   737 => x"38728407",
   738 => x"5373812a",
   739 => x"70810651",
   740 => x"5271802e",
   741 => x"85387282",
   742 => x"07537382",
   743 => x"2a708106",
   744 => x"51527180",
   745 => x"2e853872",
   746 => x"81075373",
   747 => x"832a7081",
   748 => x"06515271",
   749 => x"802e8538",
   750 => x"72880753",
   751 => x"73842a70",
   752 => x"81065152",
   753 => x"71802e85",
   754 => x"38729007",
   755 => x"5373852a",
   756 => x"70810651",
   757 => x"5271802e",
   758 => x"853872a0",
   759 => x"075372fc",
   760 => x"0c865280",
   761 => x"cbf40883",
   762 => x"38845271",
   763 => x"ec0c96e9",
   764 => x"04800b80",
   765 => x"cbf40c02",
   766 => x"90050d04",
   767 => x"71980c04",
   768 => x"ffb00880",
   769 => x"cbf40c04",
   770 => x"810bffb0",
   771 => x"0c04800b",
   772 => x"ffb00c04",
   773 => x"02f4050d",
   774 => x"99a20480",
   775 => x"cbf40881",
   776 => x"f02e0981",
   777 => x"068a3881",
   778 => x"0b80ca80",
   779 => x"0c99a204",
   780 => x"80cbf408",
   781 => x"81e02e09",
   782 => x"81068a38",
   783 => x"810b80ca",
   784 => x"840c99a2",
   785 => x"0480cbf4",
   786 => x"085280ca",
   787 => x"8408802e",
   788 => x"893880cb",
   789 => x"f4088180",
   790 => x"05527184",
   791 => x"2c728f06",
   792 => x"535380ca",
   793 => x"8008802e",
   794 => x"9a387284",
   795 => x"2980c9c0",
   796 => x"05721381",
   797 => x"712b7009",
   798 => x"73080673",
   799 => x"0c515353",
   800 => x"99960472",
   801 => x"842980c9",
   802 => x"c0057213",
   803 => x"83712b72",
   804 => x"0807720c",
   805 => x"5353800b",
   806 => x"80ca840c",
   807 => x"800b80ca",
   808 => x"800c80cc",
   809 => x"9c519aa9",
   810 => x"2d80cbf4",
   811 => x"08ff24fe",
   812 => x"ea38800b",
   813 => x"80cbf40c",
   814 => x"028c050d",
   815 => x"0402f805",
   816 => x"0d80c9c0",
   817 => x"528f5180",
   818 => x"72708405",
   819 => x"540cff11",
   820 => x"51708025",
   821 => x"f2380288",
   822 => x"050d0402",
   823 => x"f0050d75",
   824 => x"51988e2d",
   825 => x"70822cfc",
   826 => x"0680c9c0",
   827 => x"1172109e",
   828 => x"06710870",
   829 => x"722a7083",
   830 => x"0682742b",
   831 => x"70097406",
   832 => x"760c5451",
   833 => x"56575351",
   834 => x"5398882d",
   835 => x"7180cbf4",
   836 => x"0c029005",
   837 => x"0d0402fc",
   838 => x"050d7251",
   839 => x"80710c80",
   840 => x"0b84120c",
   841 => x"0284050d",
   842 => x"0402f005",
   843 => x"0d757008",
   844 => x"84120853",
   845 => x"5353ff54",
   846 => x"71712ea8",
   847 => x"38988e2d",
   848 => x"84130870",
   849 => x"84291488",
   850 => x"11700870",
   851 => x"81ff0684",
   852 => x"18088111",
   853 => x"8706841a",
   854 => x"0c535155",
   855 => x"51515198",
   856 => x"882d7154",
   857 => x"7380cbf4",
   858 => x"0c029005",
   859 => x"0d0402f8",
   860 => x"050d988e",
   861 => x"2de00870",
   862 => x"8b2a7081",
   863 => x"06515252",
   864 => x"70802ea1",
   865 => x"3880cc9c",
   866 => x"08708429",
   867 => x"80cca405",
   868 => x"7381ff06",
   869 => x"710c5151",
   870 => x"80cc9c08",
   871 => x"81118706",
   872 => x"80cc9c0c",
   873 => x"51800b80",
   874 => x"ccc40c98",
   875 => x"802d9888",
   876 => x"2d028805",
   877 => x"0d0402fc",
   878 => x"050d988e",
   879 => x"2d810b80",
   880 => x"ccc40c98",
   881 => x"882d80cc",
   882 => x"c4085170",
   883 => x"f9380284",
   884 => x"050d0402",
   885 => x"fc050d80",
   886 => x"cc9c519a",
   887 => x"962d99bd",
   888 => x"2d9aee51",
   889 => x"97fc2d02",
   890 => x"84050d04",
   891 => x"80cccc08",
   892 => x"80cbf40c",
   893 => x"0402fc05",
   894 => x"0d810b80",
   895 => x"cab40c81",
   896 => x"51858d2d",
   897 => x"0284050d",
   898 => x"0402fc05",
   899 => x"0d9c9304",
   900 => x"98942d80",
   901 => x"f65199db",
   902 => x"2d80cbf4",
   903 => x"08f23880",
   904 => x"da5199db",
   905 => x"2d80cbf4",
   906 => x"08e63880",
   907 => x"cab00851",
   908 => x"99db2d80",
   909 => x"cbf408d8",
   910 => x"3880cbf4",
   911 => x"0880cab4",
   912 => x"0c80cbf4",
   913 => x"0851858d",
   914 => x"2d028405",
   915 => x"0d0402ec",
   916 => x"050d7654",
   917 => x"8052870b",
   918 => x"881580f5",
   919 => x"2d565374",
   920 => x"72248338",
   921 => x"a0537251",
   922 => x"83842d81",
   923 => x"128b1580",
   924 => x"f52d5452",
   925 => x"727225de",
   926 => x"38029405",
   927 => x"0d0402f0",
   928 => x"050d80cc",
   929 => x"cc085481",
   930 => x"f92d800b",
   931 => x"80ccd00c",
   932 => x"7308802e",
   933 => x"81893882",
   934 => x"0b80cc88",
   935 => x"0c80ccd0",
   936 => x"088f0680",
   937 => x"cc840c73",
   938 => x"08527183",
   939 => x"2e963871",
   940 => x"83268938",
   941 => x"71812eb0",
   942 => x"389e8804",
   943 => x"71852ea0",
   944 => x"389e8804",
   945 => x"881480f5",
   946 => x"2d841508",
   947 => x"80c6a453",
   948 => x"545286a3",
   949 => x"2d718429",
   950 => x"13700852",
   951 => x"529e8c04",
   952 => x"73519cce",
   953 => x"2d9e8804",
   954 => x"80ca8808",
   955 => x"8815082c",
   956 => x"70810651",
   957 => x"5271802e",
   958 => x"883880c6",
   959 => x"a8519e85",
   960 => x"0480c6ac",
   961 => x"5186a32d",
   962 => x"84140851",
   963 => x"86a32d80",
   964 => x"ccd00881",
   965 => x"0580ccd0",
   966 => x"0c8c1454",
   967 => x"9d900402",
   968 => x"90050d04",
   969 => x"7180cccc",
   970 => x"0c9cfe2d",
   971 => x"80ccd008",
   972 => x"ff0580cc",
   973 => x"d40c0402",
   974 => x"e8050d80",
   975 => x"cccc0880",
   976 => x"ccd80857",
   977 => x"5580f651",
   978 => x"99db2d80",
   979 => x"cbf40881",
   980 => x"2a708106",
   981 => x"51527180",
   982 => x"2ea2389e",
   983 => x"e1049894",
   984 => x"2d80f651",
   985 => x"99db2d80",
   986 => x"cbf408f2",
   987 => x"3880cab4",
   988 => x"08813270",
   989 => x"80cab40c",
   990 => x"51858d2d",
   991 => x"800b80cc",
   992 => x"c80c8c51",
   993 => x"99db2d80",
   994 => x"cbf40881",
   995 => x"2a708106",
   996 => x"51527180",
   997 => x"2e80d338",
   998 => x"80ca8c08",
   999 => x"80caa008",
  1000 => x"80ca8c0c",
  1001 => x"80caa00c",
  1002 => x"80ca9008",
  1003 => x"80caa408",
  1004 => x"80ca900c",
  1005 => x"80caa40c",
  1006 => x"80ca9408",
  1007 => x"80caa808",
  1008 => x"80ca940c",
  1009 => x"80caa80c",
  1010 => x"80ca9808",
  1011 => x"80caac08",
  1012 => x"80ca980c",
  1013 => x"80caac0c",
  1014 => x"80ca9c08",
  1015 => x"80cab008",
  1016 => x"80ca9c0c",
  1017 => x"7080cab0",
  1018 => x"0c5280ca",
  1019 => x"b4088293",
  1020 => x"3880caa0",
  1021 => x"085199db",
  1022 => x"2d80cbf4",
  1023 => x"08802e8b",
  1024 => x"3880ccc8",
  1025 => x"08810780",
  1026 => x"ccc80c80",
  1027 => x"caa40851",
  1028 => x"99db2d80",
  1029 => x"cbf40880",
  1030 => x"2e8b3880",
  1031 => x"ccc80882",
  1032 => x"0780ccc8",
  1033 => x"0c80caa8",
  1034 => x"085199db",
  1035 => x"2d80cbf4",
  1036 => x"08802e8b",
  1037 => x"3880ccc8",
  1038 => x"08840780",
  1039 => x"ccc80c80",
  1040 => x"caac0851",
  1041 => x"99db2d80",
  1042 => x"cbf40880",
  1043 => x"2e8b3880",
  1044 => x"ccc80888",
  1045 => x"0780ccc8",
  1046 => x"0c80cab0",
  1047 => x"085199db",
  1048 => x"2d80cbf4",
  1049 => x"08802e8b",
  1050 => x"3880ccc8",
  1051 => x"08900780",
  1052 => x"ccc80c80",
  1053 => x"ca8c0851",
  1054 => x"99db2d80",
  1055 => x"cbf40880",
  1056 => x"2e8c3880",
  1057 => x"ccc80882",
  1058 => x"800780cc",
  1059 => x"c80c80ca",
  1060 => x"90085199",
  1061 => x"db2d80cb",
  1062 => x"f408802e",
  1063 => x"8c3880cc",
  1064 => x"c8088480",
  1065 => x"0780ccc8",
  1066 => x"0c80ca94",
  1067 => x"085199db",
  1068 => x"2d80cbf4",
  1069 => x"08802e8c",
  1070 => x"3880ccc8",
  1071 => x"08888007",
  1072 => x"80ccc80c",
  1073 => x"80ca9808",
  1074 => x"5199db2d",
  1075 => x"80cbf408",
  1076 => x"802e8c38",
  1077 => x"80ccc808",
  1078 => x"90800780",
  1079 => x"ccc80c80",
  1080 => x"ca9c0851",
  1081 => x"99db2d80",
  1082 => x"cbf40880",
  1083 => x"2e8c3880",
  1084 => x"ccc808a0",
  1085 => x"800780cc",
  1086 => x"c80c80cc",
  1087 => x"c808ed0c",
  1088 => x"a8c60481",
  1089 => x"f55199db",
  1090 => x"2d80cbf4",
  1091 => x"08812a70",
  1092 => x"81065152",
  1093 => x"71993880",
  1094 => x"caa00851",
  1095 => x"99db2d80",
  1096 => x"cbf40881",
  1097 => x"2a708106",
  1098 => x"51527180",
  1099 => x"2eb33880",
  1100 => x"ccd40852",
  1101 => x"71802e8a",
  1102 => x"38ff1280",
  1103 => x"ccd40ca2",
  1104 => x"e10480cc",
  1105 => x"d0081080",
  1106 => x"ccd00805",
  1107 => x"70842916",
  1108 => x"51528812",
  1109 => x"08802e89",
  1110 => x"38ff5188",
  1111 => x"12085271",
  1112 => x"2d81f251",
  1113 => x"99db2d80",
  1114 => x"cbf40881",
  1115 => x"2a708106",
  1116 => x"51527199",
  1117 => x"3880caa4",
  1118 => x"085199db",
  1119 => x"2d80cbf4",
  1120 => x"08812a70",
  1121 => x"81065152",
  1122 => x"71802eb4",
  1123 => x"3880ccd0",
  1124 => x"08ff1180",
  1125 => x"ccd40856",
  1126 => x"53537372",
  1127 => x"258a3881",
  1128 => x"1480ccd4",
  1129 => x"0ca3c004",
  1130 => x"72101370",
  1131 => x"84291651",
  1132 => x"52881208",
  1133 => x"802e8938",
  1134 => x"fe518812",
  1135 => x"0852712d",
  1136 => x"81fd5199",
  1137 => x"db2d80cb",
  1138 => x"f408812a",
  1139 => x"70810651",
  1140 => x"52719938",
  1141 => x"80caa808",
  1142 => x"5199db2d",
  1143 => x"80cbf408",
  1144 => x"812a7081",
  1145 => x"06515271",
  1146 => x"802eb138",
  1147 => x"80ccd408",
  1148 => x"802e8a38",
  1149 => x"800b80cc",
  1150 => x"d40ca49c",
  1151 => x"0480ccd0",
  1152 => x"081080cc",
  1153 => x"d0080570",
  1154 => x"84291651",
  1155 => x"52881208",
  1156 => x"802e8938",
  1157 => x"fd518812",
  1158 => x"0852712d",
  1159 => x"81fa5199",
  1160 => x"db2d80cb",
  1161 => x"f408812a",
  1162 => x"70810651",
  1163 => x"52719938",
  1164 => x"80caac08",
  1165 => x"5199db2d",
  1166 => x"80cbf408",
  1167 => x"812a7081",
  1168 => x"06515271",
  1169 => x"802eb138",
  1170 => x"80ccd008",
  1171 => x"ff115452",
  1172 => x"80ccd408",
  1173 => x"73258938",
  1174 => x"7280ccd4",
  1175 => x"0ca4f804",
  1176 => x"71101270",
  1177 => x"84291651",
  1178 => x"52881208",
  1179 => x"802e8938",
  1180 => x"fc518812",
  1181 => x"0852712d",
  1182 => x"80ccd408",
  1183 => x"70535473",
  1184 => x"802e8a38",
  1185 => x"8c15ff15",
  1186 => x"5555a4ff",
  1187 => x"04820b80",
  1188 => x"cc880c71",
  1189 => x"8f0680cc",
  1190 => x"840c81eb",
  1191 => x"5199db2d",
  1192 => x"80cbf408",
  1193 => x"812a7081",
  1194 => x"06515271",
  1195 => x"802ead38",
  1196 => x"7408852e",
  1197 => x"098106a4",
  1198 => x"38881580",
  1199 => x"f52dff05",
  1200 => x"52718816",
  1201 => x"81b72d71",
  1202 => x"982b5271",
  1203 => x"80258838",
  1204 => x"800b8816",
  1205 => x"81b72d74",
  1206 => x"519cce2d",
  1207 => x"81f45199",
  1208 => x"db2d80cb",
  1209 => x"f408812a",
  1210 => x"70810651",
  1211 => x"5271802e",
  1212 => x"b3387408",
  1213 => x"852e0981",
  1214 => x"06aa3888",
  1215 => x"1580f52d",
  1216 => x"81055271",
  1217 => x"881681b7",
  1218 => x"2d7181ff",
  1219 => x"068b1680",
  1220 => x"f52d5452",
  1221 => x"72722787",
  1222 => x"38728816",
  1223 => x"81b72d74",
  1224 => x"519cce2d",
  1225 => x"80da5199",
  1226 => x"db2d80cb",
  1227 => x"f408812a",
  1228 => x"70810651",
  1229 => x"52719a38",
  1230 => x"80cab008",
  1231 => x"5199db2d",
  1232 => x"80cbf408",
  1233 => x"812a7081",
  1234 => x"06515271",
  1235 => x"802e81ad",
  1236 => x"3880cccc",
  1237 => x"0880ccd4",
  1238 => x"08555373",
  1239 => x"802e8a38",
  1240 => x"8c13ff15",
  1241 => x"5553a6db",
  1242 => x"04720852",
  1243 => x"71822ea6",
  1244 => x"38718226",
  1245 => x"89387181",
  1246 => x"2eaa38a7",
  1247 => x"fd047183",
  1248 => x"2eb43871",
  1249 => x"842e0981",
  1250 => x"0680f238",
  1251 => x"88130851",
  1252 => x"9ea42da7",
  1253 => x"fd0480cc",
  1254 => x"d4085188",
  1255 => x"13085271",
  1256 => x"2da7fd04",
  1257 => x"810b8814",
  1258 => x"082b80ca",
  1259 => x"88083280",
  1260 => x"ca880ca7",
  1261 => x"d1048813",
  1262 => x"80f52d81",
  1263 => x"058b1480",
  1264 => x"f52d5354",
  1265 => x"71742483",
  1266 => x"38805473",
  1267 => x"881481b7",
  1268 => x"2d9cfe2d",
  1269 => x"a7fd0475",
  1270 => x"08802ea4",
  1271 => x"38750851",
  1272 => x"99db2d80",
  1273 => x"cbf40881",
  1274 => x"06527180",
  1275 => x"2e8c3880",
  1276 => x"ccd40851",
  1277 => x"84160852",
  1278 => x"712d8816",
  1279 => x"5675d838",
  1280 => x"8054800b",
  1281 => x"80cc880c",
  1282 => x"738f0680",
  1283 => x"cc840ca0",
  1284 => x"527380cc",
  1285 => x"d4082e09",
  1286 => x"81069938",
  1287 => x"80ccd008",
  1288 => x"ff057432",
  1289 => x"70098105",
  1290 => x"7072079f",
  1291 => x"2a917131",
  1292 => x"51515353",
  1293 => x"71518384",
  1294 => x"2d811454",
  1295 => x"8e7425c2",
  1296 => x"3880cab4",
  1297 => x"08527180",
  1298 => x"cbf40c02",
  1299 => x"98050d04",
  1300 => x"02f4050d",
  1301 => x"d45281ff",
  1302 => x"720c7108",
  1303 => x"5381ff72",
  1304 => x"0c72882b",
  1305 => x"83fe8006",
  1306 => x"72087081",
  1307 => x"ff065152",
  1308 => x"5381ff72",
  1309 => x"0c727107",
  1310 => x"882b7208",
  1311 => x"7081ff06",
  1312 => x"51525381",
  1313 => x"ff720c72",
  1314 => x"7107882b",
  1315 => x"72087081",
  1316 => x"ff067207",
  1317 => x"80cbf40c",
  1318 => x"5253028c",
  1319 => x"050d0402",
  1320 => x"f4050d74",
  1321 => x"767181ff",
  1322 => x"06d40c53",
  1323 => x"5380ccdc",
  1324 => x"08853871",
  1325 => x"892b5271",
  1326 => x"982ad40c",
  1327 => x"71902a70",
  1328 => x"81ff06d4",
  1329 => x"0c517188",
  1330 => x"2a7081ff",
  1331 => x"06d40c51",
  1332 => x"7181ff06",
  1333 => x"d40c7290",
  1334 => x"2a7081ff",
  1335 => x"06d40c51",
  1336 => x"d4087081",
  1337 => x"ff065151",
  1338 => x"82b8bf52",
  1339 => x"7081ff2e",
  1340 => x"09810694",
  1341 => x"3881ff0b",
  1342 => x"d40cd408",
  1343 => x"7081ff06",
  1344 => x"ff145451",
  1345 => x"5171e538",
  1346 => x"7080cbf4",
  1347 => x"0c028c05",
  1348 => x"0d0402fc",
  1349 => x"050d81c7",
  1350 => x"5181ff0b",
  1351 => x"d40cff11",
  1352 => x"51708025",
  1353 => x"f4380284",
  1354 => x"050d0402",
  1355 => x"f4050d81",
  1356 => x"ff0bd40c",
  1357 => x"93538052",
  1358 => x"87fc80c1",
  1359 => x"51a99f2d",
  1360 => x"80cbf408",
  1361 => x"8b3881ff",
  1362 => x"0bd40c81",
  1363 => x"53aad904",
  1364 => x"aa922dff",
  1365 => x"135372de",
  1366 => x"387280cb",
  1367 => x"f40c028c",
  1368 => x"050d0402",
  1369 => x"ec050d81",
  1370 => x"0b80ccdc",
  1371 => x"0c8454d0",
  1372 => x"08708f2a",
  1373 => x"70810651",
  1374 => x"515372f3",
  1375 => x"3872d00c",
  1376 => x"aa922d80",
  1377 => x"c6b05186",
  1378 => x"a32dd008",
  1379 => x"708f2a70",
  1380 => x"81065151",
  1381 => x"5372f338",
  1382 => x"810bd00c",
  1383 => x"b1538052",
  1384 => x"84d480c0",
  1385 => x"51a99f2d",
  1386 => x"80cbf408",
  1387 => x"812e9338",
  1388 => x"72822ebf",
  1389 => x"38ff1353",
  1390 => x"72e438ff",
  1391 => x"145473ff",
  1392 => x"ae38aa92",
  1393 => x"2d83aa52",
  1394 => x"849c80c8",
  1395 => x"51a99f2d",
  1396 => x"80cbf408",
  1397 => x"812e0981",
  1398 => x"069338a8",
  1399 => x"d02d80cb",
  1400 => x"f40883ff",
  1401 => x"ff065372",
  1402 => x"83aa2e9f",
  1403 => x"38aaab2d",
  1404 => x"ac860480",
  1405 => x"c6bc5186",
  1406 => x"a32d8053",
  1407 => x"addb0480",
  1408 => x"c6d45186",
  1409 => x"a32d8054",
  1410 => x"adac0481",
  1411 => x"ff0bd40c",
  1412 => x"b154aa92",
  1413 => x"2d8fcf53",
  1414 => x"805287fc",
  1415 => x"80f751a9",
  1416 => x"9f2d80cb",
  1417 => x"f4085580",
  1418 => x"cbf40881",
  1419 => x"2e098106",
  1420 => x"9c3881ff",
  1421 => x"0bd40c82",
  1422 => x"0a52849c",
  1423 => x"80e951a9",
  1424 => x"9f2d80cb",
  1425 => x"f408802e",
  1426 => x"8d38aa92",
  1427 => x"2dff1353",
  1428 => x"72c638ad",
  1429 => x"9f0481ff",
  1430 => x"0bd40c80",
  1431 => x"cbf40852",
  1432 => x"87fc80fa",
  1433 => x"51a99f2d",
  1434 => x"80cbf408",
  1435 => x"b23881ff",
  1436 => x"0bd40cd4",
  1437 => x"085381ff",
  1438 => x"0bd40c81",
  1439 => x"ff0bd40c",
  1440 => x"81ff0bd4",
  1441 => x"0c81ff0b",
  1442 => x"d40c7286",
  1443 => x"2a708106",
  1444 => x"76565153",
  1445 => x"72963880",
  1446 => x"cbf40854",
  1447 => x"adac0473",
  1448 => x"822efedb",
  1449 => x"38ff1454",
  1450 => x"73fee738",
  1451 => x"7380ccdc",
  1452 => x"0c738b38",
  1453 => x"815287fc",
  1454 => x"80d051a9",
  1455 => x"9f2d81ff",
  1456 => x"0bd40cd0",
  1457 => x"08708f2a",
  1458 => x"70810651",
  1459 => x"515372f3",
  1460 => x"3872d00c",
  1461 => x"81ff0bd4",
  1462 => x"0c815372",
  1463 => x"80cbf40c",
  1464 => x"0294050d",
  1465 => x"0402e805",
  1466 => x"0d785580",
  1467 => x"5681ff0b",
  1468 => x"d40cd008",
  1469 => x"708f2a70",
  1470 => x"81065151",
  1471 => x"5372f338",
  1472 => x"82810bd0",
  1473 => x"0c81ff0b",
  1474 => x"d40c7752",
  1475 => x"87fc80d1",
  1476 => x"51a99f2d",
  1477 => x"80dbc6df",
  1478 => x"5480cbf4",
  1479 => x"08802e8b",
  1480 => x"3880c6f4",
  1481 => x"5186a32d",
  1482 => x"aeff0481",
  1483 => x"ff0bd40c",
  1484 => x"d4087081",
  1485 => x"ff065153",
  1486 => x"7281fe2e",
  1487 => x"0981069e",
  1488 => x"3880ff53",
  1489 => x"a8d02d80",
  1490 => x"cbf40875",
  1491 => x"70840557",
  1492 => x"0cff1353",
  1493 => x"728025ec",
  1494 => x"388156ae",
  1495 => x"e404ff14",
  1496 => x"5473c838",
  1497 => x"81ff0bd4",
  1498 => x"0c81ff0b",
  1499 => x"d40cd008",
  1500 => x"708f2a70",
  1501 => x"81065151",
  1502 => x"5372f338",
  1503 => x"72d00c75",
  1504 => x"80cbf40c",
  1505 => x"0298050d",
  1506 => x"0402e805",
  1507 => x"0d77797b",
  1508 => x"58555580",
  1509 => x"53727625",
  1510 => x"a3387470",
  1511 => x"81055680",
  1512 => x"f52d7470",
  1513 => x"81055680",
  1514 => x"f52d5252",
  1515 => x"71712e86",
  1516 => x"388151af",
  1517 => x"be048113",
  1518 => x"53af9504",
  1519 => x"80517080",
  1520 => x"cbf40c02",
  1521 => x"98050d04",
  1522 => x"02ec050d",
  1523 => x"76557480",
  1524 => x"2e80c238",
  1525 => x"9a1580e0",
  1526 => x"2d51bddd",
  1527 => x"2d80cbf4",
  1528 => x"0880cbf4",
  1529 => x"0880d390",
  1530 => x"0c80cbf4",
  1531 => x"08545480",
  1532 => x"d2ec0880",
  1533 => x"2e9a3894",
  1534 => x"1580e02d",
  1535 => x"51bddd2d",
  1536 => x"80cbf408",
  1537 => x"902b83ff",
  1538 => x"f00a0670",
  1539 => x"75075153",
  1540 => x"7280d390",
  1541 => x"0c80d390",
  1542 => x"08537280",
  1543 => x"2e9d3880",
  1544 => x"d2e408fe",
  1545 => x"14712980",
  1546 => x"d2f80805",
  1547 => x"80d3940c",
  1548 => x"70842b80",
  1549 => x"d2f00c54",
  1550 => x"b0e90480",
  1551 => x"d2fc0880",
  1552 => x"d3900c80",
  1553 => x"d3800880",
  1554 => x"d3940c80",
  1555 => x"d2ec0880",
  1556 => x"2e8b3880",
  1557 => x"d2e40884",
  1558 => x"2b53b0e4",
  1559 => x"0480d384",
  1560 => x"08842b53",
  1561 => x"7280d2f0",
  1562 => x"0c029405",
  1563 => x"0d0402d8",
  1564 => x"050d800b",
  1565 => x"80d2ec0c",
  1566 => x"8454aae3",
  1567 => x"2d80cbf4",
  1568 => x"08802e97",
  1569 => x"3880cce0",
  1570 => x"528051ad",
  1571 => x"e52d80cb",
  1572 => x"f408802e",
  1573 => x"8638fe54",
  1574 => x"b1a304ff",
  1575 => x"14547380",
  1576 => x"24d83873",
  1577 => x"8d3880c7",
  1578 => x"845186a3",
  1579 => x"2d7355b6",
  1580 => x"f8048056",
  1581 => x"810b80d3",
  1582 => x"980c8853",
  1583 => x"80c79852",
  1584 => x"80cd9651",
  1585 => x"af892d80",
  1586 => x"cbf40876",
  1587 => x"2e098106",
  1588 => x"893880cb",
  1589 => x"f40880d3",
  1590 => x"980c8853",
  1591 => x"80c7a452",
  1592 => x"80cdb251",
  1593 => x"af892d80",
  1594 => x"cbf40889",
  1595 => x"3880cbf4",
  1596 => x"0880d398",
  1597 => x"0c80d398",
  1598 => x"08802e81",
  1599 => x"813880d0",
  1600 => x"a60b80f5",
  1601 => x"2d80d0a7",
  1602 => x"0b80f52d",
  1603 => x"71982b71",
  1604 => x"902b0780",
  1605 => x"d0a80b80",
  1606 => x"f52d7088",
  1607 => x"2b720780",
  1608 => x"d0a90b80",
  1609 => x"f52d7107",
  1610 => x"80d0de0b",
  1611 => x"80f52d80",
  1612 => x"d0df0b80",
  1613 => x"f52d7188",
  1614 => x"2b07535f",
  1615 => x"54525a56",
  1616 => x"57557381",
  1617 => x"abaa2e09",
  1618 => x"81068e38",
  1619 => x"7551bdac",
  1620 => x"2d80cbf4",
  1621 => x"0856b2e7",
  1622 => x"047382d4",
  1623 => x"d52e8838",
  1624 => x"80c7b051",
  1625 => x"b3b30480",
  1626 => x"cce05275",
  1627 => x"51ade52d",
  1628 => x"80cbf408",
  1629 => x"5580cbf4",
  1630 => x"08802e83",
  1631 => x"fb388853",
  1632 => x"80c7a452",
  1633 => x"80cdb251",
  1634 => x"af892d80",
  1635 => x"cbf4088a",
  1636 => x"38810b80",
  1637 => x"d2ec0cb3",
  1638 => x"b9048853",
  1639 => x"80c79852",
  1640 => x"80cd9651",
  1641 => x"af892d80",
  1642 => x"cbf40880",
  1643 => x"2e8b3880",
  1644 => x"c7c45186",
  1645 => x"a32db498",
  1646 => x"0480d0de",
  1647 => x"0b80f52d",
  1648 => x"547380d5",
  1649 => x"2e098106",
  1650 => x"80ce3880",
  1651 => x"d0df0b80",
  1652 => x"f52d5473",
  1653 => x"81aa2e09",
  1654 => x"8106bd38",
  1655 => x"800b80cc",
  1656 => x"e00b80f5",
  1657 => x"2d565474",
  1658 => x"81e92e83",
  1659 => x"38815474",
  1660 => x"81eb2e8c",
  1661 => x"38805573",
  1662 => x"752e0981",
  1663 => x"0682f938",
  1664 => x"80cceb0b",
  1665 => x"80f52d55",
  1666 => x"748e3880",
  1667 => x"ccec0b80",
  1668 => x"f52d5473",
  1669 => x"822e8638",
  1670 => x"8055b6f8",
  1671 => x"0480cced",
  1672 => x"0b80f52d",
  1673 => x"7080d2e4",
  1674 => x"0cff0580",
  1675 => x"d2e80c80",
  1676 => x"ccee0b80",
  1677 => x"f52d80cc",
  1678 => x"ef0b80f5",
  1679 => x"2d587605",
  1680 => x"77828029",
  1681 => x"057080d2",
  1682 => x"f40c80cc",
  1683 => x"f00b80f5",
  1684 => x"2d7080d3",
  1685 => x"880c80d2",
  1686 => x"ec085957",
  1687 => x"5876802e",
  1688 => x"81b73888",
  1689 => x"5380c7a4",
  1690 => x"5280cdb2",
  1691 => x"51af892d",
  1692 => x"80cbf408",
  1693 => x"82823880",
  1694 => x"d2e40870",
  1695 => x"842b80d2",
  1696 => x"f00c7080",
  1697 => x"d3840c80",
  1698 => x"cd850b80",
  1699 => x"f52d80cd",
  1700 => x"840b80f5",
  1701 => x"2d718280",
  1702 => x"290580cd",
  1703 => x"860b80f5",
  1704 => x"2d708480",
  1705 => x"80291280",
  1706 => x"cd870b80",
  1707 => x"f52d7081",
  1708 => x"800a2912",
  1709 => x"7080d38c",
  1710 => x"0c80d388",
  1711 => x"08712980",
  1712 => x"d2f40805",
  1713 => x"7080d2f8",
  1714 => x"0c80cd8d",
  1715 => x"0b80f52d",
  1716 => x"80cd8c0b",
  1717 => x"80f52d71",
  1718 => x"82802905",
  1719 => x"80cd8e0b",
  1720 => x"80f52d70",
  1721 => x"84808029",
  1722 => x"1280cd8f",
  1723 => x"0b80f52d",
  1724 => x"70982b81",
  1725 => x"f00a0672",
  1726 => x"057080d2",
  1727 => x"fc0cfe11",
  1728 => x"7e297705",
  1729 => x"80d3800c",
  1730 => x"52595243",
  1731 => x"545e5152",
  1732 => x"59525d57",
  1733 => x"5957b6f1",
  1734 => x"0480ccf2",
  1735 => x"0b80f52d",
  1736 => x"80ccf10b",
  1737 => x"80f52d71",
  1738 => x"82802905",
  1739 => x"7080d2f0",
  1740 => x"0c70a029",
  1741 => x"83ff0570",
  1742 => x"892a7080",
  1743 => x"d3840c80",
  1744 => x"ccf70b80",
  1745 => x"f52d80cc",
  1746 => x"f60b80f5",
  1747 => x"2d718280",
  1748 => x"29057080",
  1749 => x"d38c0c7b",
  1750 => x"71291e70",
  1751 => x"80d3800c",
  1752 => x"7d80d2fc",
  1753 => x"0c730580",
  1754 => x"d2f80c55",
  1755 => x"5e515155",
  1756 => x"558051af",
  1757 => x"c82d8155",
  1758 => x"7480cbf4",
  1759 => x"0c02a805",
  1760 => x"0d0402ec",
  1761 => x"050d7670",
  1762 => x"872c7180",
  1763 => x"ff065556",
  1764 => x"5480d2ec",
  1765 => x"088a3873",
  1766 => x"882c7481",
  1767 => x"ff065455",
  1768 => x"80cce052",
  1769 => x"80d2f408",
  1770 => x"1551ade5",
  1771 => x"2d80cbf4",
  1772 => x"085480cb",
  1773 => x"f408802e",
  1774 => x"b83880d2",
  1775 => x"ec08802e",
  1776 => x"9a387284",
  1777 => x"2980cce0",
  1778 => x"05700852",
  1779 => x"53bdac2d",
  1780 => x"80cbf408",
  1781 => x"f00a0653",
  1782 => x"b7ef0472",
  1783 => x"1080cce0",
  1784 => x"057080e0",
  1785 => x"2d5253bd",
  1786 => x"dd2d80cb",
  1787 => x"f4085372",
  1788 => x"547380cb",
  1789 => x"f40c0294",
  1790 => x"050d0402",
  1791 => x"e0050d79",
  1792 => x"70842c80",
  1793 => x"d3940805",
  1794 => x"718f0652",
  1795 => x"5553728a",
  1796 => x"3880cce0",
  1797 => x"527351ad",
  1798 => x"e52d72a0",
  1799 => x"2980cce0",
  1800 => x"05548074",
  1801 => x"80f52d56",
  1802 => x"5374732e",
  1803 => x"83388153",
  1804 => x"7481e52e",
  1805 => x"81f43881",
  1806 => x"70740654",
  1807 => x"5872802e",
  1808 => x"81e8388b",
  1809 => x"1480f52d",
  1810 => x"70832a79",
  1811 => x"06585676",
  1812 => x"9b3880ca",
  1813 => x"b8085372",
  1814 => x"89387280",
  1815 => x"d0e00b81",
  1816 => x"b72d7680",
  1817 => x"cab80c73",
  1818 => x"53baac04",
  1819 => x"758f2e09",
  1820 => x"810681b6",
  1821 => x"38749f06",
  1822 => x"8d2980d0",
  1823 => x"d3115153",
  1824 => x"811480f5",
  1825 => x"2d737081",
  1826 => x"055581b7",
  1827 => x"2d831480",
  1828 => x"f52d7370",
  1829 => x"81055581",
  1830 => x"b72d8514",
  1831 => x"80f52d73",
  1832 => x"70810555",
  1833 => x"81b72d87",
  1834 => x"1480f52d",
  1835 => x"73708105",
  1836 => x"5581b72d",
  1837 => x"891480f5",
  1838 => x"2d737081",
  1839 => x"055581b7",
  1840 => x"2d8e1480",
  1841 => x"f52d7370",
  1842 => x"81055581",
  1843 => x"b72d9014",
  1844 => x"80f52d73",
  1845 => x"70810555",
  1846 => x"81b72d92",
  1847 => x"1480f52d",
  1848 => x"73708105",
  1849 => x"5581b72d",
  1850 => x"941480f5",
  1851 => x"2d737081",
  1852 => x"055581b7",
  1853 => x"2d961480",
  1854 => x"f52d7370",
  1855 => x"81055581",
  1856 => x"b72d9814",
  1857 => x"80f52d73",
  1858 => x"70810555",
  1859 => x"81b72d9c",
  1860 => x"1480f52d",
  1861 => x"73708105",
  1862 => x"5581b72d",
  1863 => x"9e1480f5",
  1864 => x"2d7381b7",
  1865 => x"2d7780ca",
  1866 => x"b80c8053",
  1867 => x"7280cbf4",
  1868 => x"0c02a005",
  1869 => x"0d0402cc",
  1870 => x"050d7e60",
  1871 => x"5e5a800b",
  1872 => x"80d39008",
  1873 => x"80d39408",
  1874 => x"595c5680",
  1875 => x"5880d2f0",
  1876 => x"08782e81",
  1877 => x"b838778f",
  1878 => x"06a01757",
  1879 => x"54739138",
  1880 => x"80cce052",
  1881 => x"76518117",
  1882 => x"57ade52d",
  1883 => x"80cce056",
  1884 => x"807680f5",
  1885 => x"2d565474",
  1886 => x"742e8338",
  1887 => x"81547481",
  1888 => x"e52e80fd",
  1889 => x"38817075",
  1890 => x"06555c73",
  1891 => x"802e80f1",
  1892 => x"388b1680",
  1893 => x"f52d9806",
  1894 => x"597880e5",
  1895 => x"388b537c",
  1896 => x"527551af",
  1897 => x"892d80cb",
  1898 => x"f40880d5",
  1899 => x"389c1608",
  1900 => x"51bdac2d",
  1901 => x"80cbf408",
  1902 => x"841b0c9a",
  1903 => x"1680e02d",
  1904 => x"51bddd2d",
  1905 => x"80cbf408",
  1906 => x"80cbf408",
  1907 => x"881c0c80",
  1908 => x"cbf40855",
  1909 => x"5580d2ec",
  1910 => x"08802e99",
  1911 => x"38941680",
  1912 => x"e02d51bd",
  1913 => x"dd2d80cb",
  1914 => x"f408902b",
  1915 => x"83fff00a",
  1916 => x"06701651",
  1917 => x"5473881b",
  1918 => x"0c787a0c",
  1919 => x"7b54bcc9",
  1920 => x"04811858",
  1921 => x"80d2f008",
  1922 => x"7826feca",
  1923 => x"3880d2ec",
  1924 => x"08802eb3",
  1925 => x"387a51b7",
  1926 => x"822d80cb",
  1927 => x"f40880cb",
  1928 => x"f40880ff",
  1929 => x"fffff806",
  1930 => x"555b7380",
  1931 => x"fffffff8",
  1932 => x"2e953880",
  1933 => x"cbf408fe",
  1934 => x"0580d2e4",
  1935 => x"082980d2",
  1936 => x"f8080557",
  1937 => x"bacb0480",
  1938 => x"547380cb",
  1939 => x"f40c02b4",
  1940 => x"050d0402",
  1941 => x"f4050d74",
  1942 => x"70088105",
  1943 => x"710c7008",
  1944 => x"80d2e808",
  1945 => x"06535371",
  1946 => x"8f388813",
  1947 => x"0851b782",
  1948 => x"2d80cbf4",
  1949 => x"0888140c",
  1950 => x"810b80cb",
  1951 => x"f40c028c",
  1952 => x"050d0402",
  1953 => x"f0050d75",
  1954 => x"881108fe",
  1955 => x"0580d2e4",
  1956 => x"082980d2",
  1957 => x"f8081172",
  1958 => x"0880d2e8",
  1959 => x"08060579",
  1960 => x"55535454",
  1961 => x"ade52d02",
  1962 => x"90050d04",
  1963 => x"02f4050d",
  1964 => x"7470882a",
  1965 => x"83fe8006",
  1966 => x"7072982a",
  1967 => x"0772882b",
  1968 => x"87fc8080",
  1969 => x"0673982b",
  1970 => x"81f00a06",
  1971 => x"71730707",
  1972 => x"80cbf40c",
  1973 => x"56515351",
  1974 => x"028c050d",
  1975 => x"0402f805",
  1976 => x"0d028e05",
  1977 => x"80f52d74",
  1978 => x"882b0770",
  1979 => x"83ffff06",
  1980 => x"80cbf40c",
  1981 => x"51028805",
  1982 => x"0d0402f4",
  1983 => x"050d7476",
  1984 => x"78535452",
  1985 => x"80712597",
  1986 => x"38727081",
  1987 => x"055480f5",
  1988 => x"2d727081",
  1989 => x"055481b7",
  1990 => x"2dff1151",
  1991 => x"70eb3880",
  1992 => x"7281b72d",
  1993 => x"028c050d",
  1994 => x"0402e805",
  1995 => x"0d775680",
  1996 => x"70565473",
  1997 => x"7624b638",
  1998 => x"80d2f008",
  1999 => x"742eae38",
  2000 => x"7351b7fb",
  2001 => x"2d80cbf4",
  2002 => x"0880cbf4",
  2003 => x"08098105",
  2004 => x"7080cbf4",
  2005 => x"08079f2a",
  2006 => x"77058117",
  2007 => x"57575353",
  2008 => x"74762489",
  2009 => x"3880d2f0",
  2010 => x"087426d4",
  2011 => x"387280cb",
  2012 => x"f40c0298",
  2013 => x"050d0402",
  2014 => x"f0050d80",
  2015 => x"cbf00816",
  2016 => x"51bea92d",
  2017 => x"80cbf408",
  2018 => x"802e9f38",
  2019 => x"8b5380cb",
  2020 => x"f4085280",
  2021 => x"d0e051bd",
  2022 => x"fa2d80d3",
  2023 => x"9c085473",
  2024 => x"802e8738",
  2025 => x"80d0e051",
  2026 => x"732d0290",
  2027 => x"050d0402",
  2028 => x"dc050d80",
  2029 => x"705a5574",
  2030 => x"80cbf008",
  2031 => x"25b43880",
  2032 => x"d2f00875",
  2033 => x"2eac3878",
  2034 => x"51b7fb2d",
  2035 => x"80cbf408",
  2036 => x"09810570",
  2037 => x"80cbf408",
  2038 => x"079f2a76",
  2039 => x"05811b5b",
  2040 => x"56547480",
  2041 => x"cbf00825",
  2042 => x"893880d2",
  2043 => x"f0087926",
  2044 => x"d6388055",
  2045 => x"7880d2f0",
  2046 => x"082781e0",
  2047 => x"387851b7",
  2048 => x"fb2d80cb",
  2049 => x"f408802e",
  2050 => x"81b23880",
  2051 => x"cbf4088b",
  2052 => x"0580f52d",
  2053 => x"70842a70",
  2054 => x"81067710",
  2055 => x"78842b80",
  2056 => x"d0e00b80",
  2057 => x"f52d5c5c",
  2058 => x"53515556",
  2059 => x"73802e80",
  2060 => x"ce387416",
  2061 => x"822b80c2",
  2062 => x"800b80ca",
  2063 => x"c4120c54",
  2064 => x"77753110",
  2065 => x"80d3a011",
  2066 => x"55569074",
  2067 => x"70810556",
  2068 => x"81b72da0",
  2069 => x"7481b72d",
  2070 => x"7681ff06",
  2071 => x"81165854",
  2072 => x"73802e8b",
  2073 => x"389c5380",
  2074 => x"d0e05280",
  2075 => x"c0f6048b",
  2076 => x"5380cbf4",
  2077 => x"085280d3",
  2078 => x"a2165180",
  2079 => x"c1b30474",
  2080 => x"16822bbe",
  2081 => x"f70b80ca",
  2082 => x"c4120c54",
  2083 => x"7681ff06",
  2084 => x"81165854",
  2085 => x"73802e8b",
  2086 => x"389c5380",
  2087 => x"d0e05280",
  2088 => x"c1aa048b",
  2089 => x"5380cbf4",
  2090 => x"08527775",
  2091 => x"311080d3",
  2092 => x"a0055176",
  2093 => x"55bdfa2d",
  2094 => x"80c1d104",
  2095 => x"74902975",
  2096 => x"31701080",
  2097 => x"d3a00551",
  2098 => x"5480cbf4",
  2099 => x"087481b7",
  2100 => x"2d811959",
  2101 => x"748b24a3",
  2102 => x"38bff404",
  2103 => x"74902975",
  2104 => x"31701080",
  2105 => x"d3a0058c",
  2106 => x"77315751",
  2107 => x"54807481",
  2108 => x"b72d9e14",
  2109 => x"ff165654",
  2110 => x"74f33802",
  2111 => x"a4050d04",
  2112 => x"02fc050d",
  2113 => x"80cbf008",
  2114 => x"1351bea9",
  2115 => x"2d80cbf4",
  2116 => x"08802e89",
  2117 => x"3880cbf4",
  2118 => x"0851afc8",
  2119 => x"2d800b80",
  2120 => x"cbf00cbf",
  2121 => x"af2d9cfe",
  2122 => x"2d028405",
  2123 => x"0d0402fc",
  2124 => x"050d7251",
  2125 => x"70fd2eb2",
  2126 => x"3870fd24",
  2127 => x"8b3870fc",
  2128 => x"2e80d038",
  2129 => x"80c39d04",
  2130 => x"70fe2eb9",
  2131 => x"3870ff2e",
  2132 => x"09810680",
  2133 => x"c83880cb",
  2134 => x"f0085170",
  2135 => x"802ebe38",
  2136 => x"ff1180cb",
  2137 => x"f00c80c3",
  2138 => x"9d0480cb",
  2139 => x"f008f405",
  2140 => x"7080cbf0",
  2141 => x"0c517080",
  2142 => x"25a33880",
  2143 => x"0b80cbf0",
  2144 => x"0c80c39d",
  2145 => x"0480cbf0",
  2146 => x"08810580",
  2147 => x"cbf00c80",
  2148 => x"c39d0480",
  2149 => x"cbf0088c",
  2150 => x"0580cbf0",
  2151 => x"0cbfaf2d",
  2152 => x"9cfe2d02",
  2153 => x"84050d04",
  2154 => x"02fc050d",
  2155 => x"800b80cb",
  2156 => x"f00cbfaf",
  2157 => x"2d9bec2d",
  2158 => x"80cbf408",
  2159 => x"80cbe00c",
  2160 => x"80cabc51",
  2161 => x"9ea42d02",
  2162 => x"84050d04",
  2163 => x"7180d39c",
  2164 => x"0c040000",
  2165 => x"00ffffff",
  2166 => x"ff00ffff",
  2167 => x"ffff00ff",
  2168 => x"ffffff00",
  2169 => x"436f6e74",
  2170 => x"696e7565",
  2171 => x"00000000",
  2172 => x"52657365",
  2173 => x"74000000",
  2174 => x"446f7562",
  2175 => x"6c65204f",
  2176 => x"53442077",
  2177 => x"696e646f",
  2178 => x"77000000",
  2179 => x"4c6f6164",
  2180 => x"20546170",
  2181 => x"6520282e",
  2182 => x"702c202e",
  2183 => x"38312920",
  2184 => x"10000000",
  2185 => x"45786974",
  2186 => x"00000000",
  2187 => x"524f4d20",
  2188 => x"6c6f6164",
  2189 => x"696e6720",
  2190 => x"6661696c",
  2191 => x"65640000",
  2192 => x"4f4b0000",
  2193 => x"54617065",
  2194 => x"2066696c",
  2195 => x"65204c6f",
  2196 => x"61646564",
  2197 => x"2e000000",
  2198 => x"54797065",
  2199 => x"204c4f41",
  2200 => x"44202222",
  2201 => x"202b2045",
  2202 => x"4e544552",
  2203 => x"206f6e20",
  2204 => x"5a583831",
  2205 => x"00000000",
  2206 => x"5468656e",
  2207 => x"20707265",
  2208 => x"73732050",
  2209 => x"6c617920",
  2210 => x"616e6420",
  2211 => x"77616974",
  2212 => x"00000000",
  2213 => x"54686572",
  2214 => x"65206973",
  2215 => x"206e6f20",
  2216 => x"696d6167",
  2217 => x"65207768",
  2218 => x"656e206c",
  2219 => x"6f616469",
  2220 => x"6e670000",
  2221 => x"54617065",
  2222 => x"204b6579",
  2223 => x"733a0000",
  2224 => x"20202d20",
  2225 => x"46353a20",
  2226 => x"506c6179",
  2227 => x"2f506175",
  2228 => x"73650000",
  2229 => x"20202d20",
  2230 => x"46363a20",
  2231 => x"53746f70",
  2232 => x"20746865",
  2233 => x"20746170",
  2234 => x"65000000",
  2235 => x"20202d20",
  2236 => x"46373a20",
  2237 => x"456a6563",
  2238 => x"74202d28",
  2239 => x"52657365",
  2240 => x"74732074",
  2241 => x"61706529",
  2242 => x"00000000",
  2243 => x"496e6974",
  2244 => x"69616c69",
  2245 => x"7a696e67",
  2246 => x"20534420",
  2247 => x"63617264",
  2248 => x"0a000000",
  2249 => x"16200000",
  2250 => x"14200000",
  2251 => x"15200000",
  2252 => x"53442069",
  2253 => x"6e69742e",
  2254 => x"2e2e0a00",
  2255 => x"53442063",
  2256 => x"61726420",
  2257 => x"72657365",
  2258 => x"74206661",
  2259 => x"696c6564",
  2260 => x"210a0000",
  2261 => x"53444843",
  2262 => x"20657272",
  2263 => x"6f72210a",
  2264 => x"00000000",
  2265 => x"57726974",
  2266 => x"65206661",
  2267 => x"696c6564",
  2268 => x"0a000000",
  2269 => x"52656164",
  2270 => x"20666169",
  2271 => x"6c65640a",
  2272 => x"00000000",
  2273 => x"43617264",
  2274 => x"20696e69",
  2275 => x"74206661",
  2276 => x"696c6564",
  2277 => x"0a000000",
  2278 => x"46415431",
  2279 => x"36202020",
  2280 => x"00000000",
  2281 => x"46415433",
  2282 => x"32202020",
  2283 => x"00000000",
  2284 => x"4e6f2070",
  2285 => x"61727469",
  2286 => x"74696f6e",
  2287 => x"20736967",
  2288 => x"0a000000",
  2289 => x"42616420",
  2290 => x"70617274",
  2291 => x"0a000000",
  2292 => x"4261636b",
  2293 => x"00000000",
  2294 => x"00000002",
  2295 => x"00000002",
  2296 => x"000021f0",
  2297 => x"0000035d",
  2298 => x"00000001",
  2299 => x"000021f8",
  2300 => x"00000005",
  2301 => x"00000002",
  2302 => x"0000220c",
  2303 => x"000021a8",
  2304 => x"00000002",
  2305 => x"00002224",
  2306 => x"00000e09",
  2307 => x"00000000",
  2308 => x"00000000",
  2309 => x"00000000",
  2310 => x"00000004",
  2311 => x"0000222c",
  2312 => x"00002418",
  2313 => x"00000004",
  2314 => x"00002240",
  2315 => x"000023dc",
  2316 => x"00000000",
  2317 => x"00000000",
  2318 => x"00000000",
  2319 => x"00000004",
  2320 => x"00002244",
  2321 => x"0000243c",
  2322 => x"00000004",
  2323 => x"00002258",
  2324 => x"0000243c",
  2325 => x"00000004",
  2326 => x"00002278",
  2327 => x"0000243c",
  2328 => x"00000004",
  2329 => x"00002294",
  2330 => x"0000243c",
  2331 => x"00000004",
  2332 => x"000022b4",
  2333 => x"0000243c",
  2334 => x"00000004",
  2335 => x"000022c0",
  2336 => x"0000243c",
  2337 => x"00000004",
  2338 => x"000022d4",
  2339 => x"0000243c",
  2340 => x"00000004",
  2341 => x"000022ec",
  2342 => x"0000243c",
  2343 => x"00000004",
  2344 => x"00002360",
  2345 => x"0000243c",
  2346 => x"00000004",
  2347 => x"000021e4",
  2348 => x"000023dc",
  2349 => x"00000000",
  2350 => x"00000000",
  2351 => x"00000000",
  2352 => x"00000000",
  2353 => x"00000000",
  2354 => x"00000000",
  2355 => x"00000000",
  2356 => x"00000000",
  2357 => x"00000000",
  2358 => x"00000000",
  2359 => x"00000000",
  2360 => x"00000000",
  2361 => x"00000000",
  2362 => x"00000000",
  2363 => x"00000000",
  2364 => x"00000000",
  2365 => x"00000000",
  2366 => x"00000000",
  2367 => x"00000000",
  2368 => x"00000000",
  2369 => x"00000000",
  2370 => x"00000006",
  2371 => x"00000043",
  2372 => x"00000042",
  2373 => x"0000003b",
  2374 => x"0000004b",
  2375 => x"00000033",
  2376 => x"00000003",
  2377 => x"0000000b",
  2378 => x"00000083",
  2379 => x"00000023",
  2380 => x"0000002b",
  2381 => x"00000000",
  2382 => x"00000000",
  2383 => x"00000002",
  2384 => x"000029a0",
  2385 => x"00001f77",
  2386 => x"00000002",
  2387 => x"000029be",
  2388 => x"00001f77",
  2389 => x"00000002",
  2390 => x"000029dc",
  2391 => x"00001f77",
  2392 => x"00000002",
  2393 => x"000029fa",
  2394 => x"00001f77",
  2395 => x"00000002",
  2396 => x"00002a18",
  2397 => x"00001f77",
  2398 => x"00000002",
  2399 => x"00002a36",
  2400 => x"00001f77",
  2401 => x"00000002",
  2402 => x"00002a54",
  2403 => x"00001f77",
  2404 => x"00000002",
  2405 => x"00002a72",
  2406 => x"00001f77",
  2407 => x"00000002",
  2408 => x"00002a90",
  2409 => x"00001f77",
  2410 => x"00000002",
  2411 => x"00002aae",
  2412 => x"00001f77",
  2413 => x"00000002",
  2414 => x"00002acc",
  2415 => x"00001f77",
  2416 => x"00000002",
  2417 => x"00002aea",
  2418 => x"00001f77",
  2419 => x"00000002",
  2420 => x"00002b08",
  2421 => x"00001f77",
  2422 => x"00000004",
  2423 => x"000023d0",
  2424 => x"00000000",
  2425 => x"00000000",
  2426 => x"00000000",
  2427 => x"0000212e",
  2428 => x"00000000",
	others => x"00000000"
);

begin

process (clk)
begin
	if (clk'event and clk = '1') then
		if (from_zpu.memAWriteEnable = '1') and (from_zpu.memBWriteEnable = '1') and (from_zpu.memAAddr=from_zpu.memBAddr) and (from_zpu.memAWrite/=from_zpu.memBWrite) then
			report "write collision" severity failure;
		end if;
	
		if (from_zpu.memAWriteEnable = '1') then
			ram(to_integer(unsigned(from_zpu.memAAddr(maxAddrBitBRAM downto 2)))) := from_zpu.memAWrite;
			to_zpu.memARead <= from_zpu.memAWrite;
		else
			to_zpu.memARead <= ram(to_integer(unsigned(from_zpu.memAAddr(maxAddrBitBRAM downto 2))));
		end if;
	end if;
end process;

process (clk)
begin
	if (clk'event and clk = '1') then
		if (from_zpu.memBWriteEnable = '1') then
			ram(to_integer(unsigned(from_zpu.memBAddr(maxAddrBitBRAM downto 2)))) := from_zpu.memBWrite;
			to_zpu.memBRead <= from_zpu.memBWrite;
		else
			to_zpu.memBRead <= ram(to_integer(unsigned(from_zpu.memBAddr(maxAddrBitBRAM downto 2))));
		end if;
	end if;
end process;


end arch;

