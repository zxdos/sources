-- ZPU
--
-- Copyright 2004-2008 oharboe - �yvind Harboe - oyvind.harboe@zylin.com
-- Modified by Alastair M. Robinson for the ZPUFlex project.
--
-- The FreeBSD license
-- 
-- Redistribution and use in source and binary forms, with or without
-- modification, are permitted provided that the following conditions
-- are met:
-- 
-- 1. Redistributions of source code must retain the above copyright
--    notice, this list of conditions and the following disclaimer.
-- 2. Redistributions in binary form must reproduce the above
--    copyright notice, this list of conditions and the following
--    disclaimer in the documentation and/or other materials
--    provided with the distribution.
-- 
-- THIS SOFTWARE IS PROVIDED BY THE ZPU PROJECT ``AS IS'' AND ANY
-- EXPRESS OR IMPLIED WARRANTIES, INCLUDING, BUT NOT LIMITED TO,
-- THE IMPLIED WARRANTIES OF MERCHANTABILITY AND FITNESS FOR A
-- PARTICULAR PURPOSE ARE DISCLAIMED. IN NO EVENT SHALL THE
-- ZPU PROJECT OR CONTRIBUTORS BE LIABLE FOR ANY DIRECT,
-- INDIRECT, INCIDENTAL, SPECIAL, EXEMPLARY, OR CONSEQUENTIAL DAMAGES
-- (INCLUDING, BUT NOT LIMITED TO, PROCUREMENT OF SUBSTITUTE GOODS
-- OR SERVICES; LOSS OF USE, DATA, OR PROFITS; OR BUSINESS INTERRUPTION)
-- HOWEVER CAUSED AND ON ANY THEORY OF LIABILITY, WHETHER IN CONTRACT,
-- STRICT LIABILITY, OR TORT (INCLUDING NEGLIGENCE OR OTHERWISE)
-- ARISING IN ANY WAY OUT OF THE USE OF THIS SOFTWARE, EVEN IF
-- ADVISED OF THE POSSIBILITY OF SUCH DAMAGE.
-- 
-- The views and conclusions contained in the software and documentation
-- are those of the authors and should not be interpreted as representing
-- official policies, either expressed or implied, of the ZPU Project.

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;


library work;
use work.zpupkg.all;

entity CtrlROM_ROM is
generic
	(
		maxAddrBitBRAM : integer := maxAddrBitBRAMLimit -- Specify your actual ROM size to save LEs and unnecessary block RAM usage.
	);
port (
	clk : in std_logic;
	areset : in std_logic := '0';
	from_zpu : in ZPU_ToROM;
	to_zpu : out ZPU_FromROM
);
end CtrlROM_ROM;

architecture arch of CtrlROM_ROM is

type ram_type is array(natural range 0 to ((2**(maxAddrBitBRAM+1))/4)-1) of std_logic_vector(wordSize-1 downto 0);

shared variable ram : ram_type :=
(
     0 => x"0b0b0b0b",
     1 => x"8c0b0b0b",
     2 => x"0b81e004",
     3 => x"0b0b0b0b",
     4 => x"8c04ff0d",
     5 => x"80040400",
     6 => x"00000016",
     7 => x"00000000",
     8 => x"0b0b0baa",
     9 => x"e4080b0b",
    10 => x"0baae808",
    11 => x"0b0b0baa",
    12 => x"ec080b0b",
    13 => x"0b0b9808",
    14 => x"2d0b0b0b",
    15 => x"aaec0c0b",
    16 => x"0b0baae8",
    17 => x"0c0b0b0b",
    18 => x"aae40c04",
    19 => x"00000000",
    20 => x"00000000",
    21 => x"00000000",
    22 => x"00000000",
    23 => x"00000000",
    24 => x"71fd0608",
    25 => x"72830609",
    26 => x"81058205",
    27 => x"832b2a83",
    28 => x"ffff0652",
    29 => x"0471fc06",
    30 => x"08728306",
    31 => x"09810583",
    32 => x"05101010",
    33 => x"2a81ff06",
    34 => x"520471fd",
    35 => x"060883ff",
    36 => x"ff738306",
    37 => x"09810582",
    38 => x"05832b2b",
    39 => x"09067383",
    40 => x"ffff0673",
    41 => x"83060981",
    42 => x"05820583",
    43 => x"2b0b2b07",
    44 => x"72fc060c",
    45 => x"51510471",
    46 => x"fc06080b",
    47 => x"0b0ba580",
    48 => x"73830610",
    49 => x"10050806",
    50 => x"7381ff06",
    51 => x"73830609",
    52 => x"81058305",
    53 => x"1010102b",
    54 => x"0772fc06",
    55 => x"0c515104",
    56 => x"aae470af",
    57 => x"fc278b38",
    58 => x"80717084",
    59 => x"05530c81",
    60 => x"e2048c51",
    61 => x"85e80402",
    62 => x"fc050df8",
    63 => x"80518f0b",
    64 => x"aaf40c9f",
    65 => x"0baaf80c",
    66 => x"a0717081",
    67 => x"055334aa",
    68 => x"f808ff05",
    69 => x"aaf80caa",
    70 => x"f8088025",
    71 => x"eb38aaf4",
    72 => x"08ff05aa",
    73 => x"f40caaf4",
    74 => x"088025d7",
    75 => x"38800baa",
    76 => x"f80c800b",
    77 => x"aaf40c02",
    78 => x"84050d04",
    79 => x"02f0050d",
    80 => x"f88053f8",
    81 => x"a05483bf",
    82 => x"52737081",
    83 => x"05553351",
    84 => x"70737081",
    85 => x"055534ff",
    86 => x"12527180",
    87 => x"25eb38fb",
    88 => x"c0539f52",
    89 => x"a0737081",
    90 => x"055534ff",
    91 => x"12527180",
    92 => x"25f23802",
    93 => x"90050d04",
    94 => x"02f4050d",
    95 => x"74538e0b",
    96 => x"aaf40825",
    97 => x"8f3882bc",
    98 => x"2daaf408",
    99 => x"ff05aaf4",
   100 => x"0c82fe04",
   101 => x"aaf408aa",
   102 => x"f8085351",
   103 => x"728a2e09",
   104 => x"8106b738",
   105 => x"7151719f",
   106 => x"24a038aa",
   107 => x"f408a029",
   108 => x"11f88011",
   109 => x"5151a071",
   110 => x"34aaf808",
   111 => x"8105aaf8",
   112 => x"0caaf808",
   113 => x"519f7125",
   114 => x"e238800b",
   115 => x"aaf80caa",
   116 => x"f4088105",
   117 => x"aaf40c83",
   118 => x"ee0470a0",
   119 => x"2912f880",
   120 => x"11515172",
   121 => x"7134aaf8",
   122 => x"088105aa",
   123 => x"f80caaf8",
   124 => x"08a02e09",
   125 => x"81068e38",
   126 => x"800baaf8",
   127 => x"0caaf408",
   128 => x"8105aaf4",
   129 => x"0c028c05",
   130 => x"0d0402ec",
   131 => x"050d800b",
   132 => x"aafc0cf6",
   133 => x"8c08f690",
   134 => x"0871882c",
   135 => x"565481ff",
   136 => x"06527372",
   137 => x"25883871",
   138 => x"54820baa",
   139 => x"fc0c7288",
   140 => x"2c7381ff",
   141 => x"06545574",
   142 => x"73258b38",
   143 => x"72aafc08",
   144 => x"8407aafc",
   145 => x"0c557384",
   146 => x"2b86a071",
   147 => x"25837131",
   148 => x"700b0b0b",
   149 => x"a8b80c81",
   150 => x"712bff05",
   151 => x"f6880cfc",
   152 => x"08fea414",
   153 => x"ff132c79",
   154 => x"8829fed0",
   155 => x"0570812c",
   156 => x"aafc0852",
   157 => x"59535155",
   158 => x"51525476",
   159 => x"802e8538",
   160 => x"70810751",
   161 => x"70f6940c",
   162 => x"71098105",
   163 => x"f6800c72",
   164 => x"098105f6",
   165 => x"840c0294",
   166 => x"050d0402",
   167 => x"f4050d74",
   168 => x"53727081",
   169 => x"055480f5",
   170 => x"2d527180",
   171 => x"2e893871",
   172 => x"5182f82d",
   173 => x"85a10481",
   174 => x"0baae40c",
   175 => x"028c050d",
   176 => x"0402fc05",
   177 => x"0d818080",
   178 => x"51c01151",
   179 => x"70fb3802",
   180 => x"84050d04",
   181 => x"02fc050d",
   182 => x"ec518371",
   183 => x"0c85c12d",
   184 => x"82710c02",
   185 => x"84050d04",
   186 => x"02f0050d",
   187 => x"805185d4",
   188 => x"2d840bec",
   189 => x"0c8b982d",
   190 => x"87e72d81",
   191 => x"f72d8352",
   192 => x"8afd2d81",
   193 => x"51848a2d",
   194 => x"ff125271",
   195 => x"8025f138",
   196 => x"840bec0c",
   197 => x"a6f45185",
   198 => x"9b2d9eef",
   199 => x"2daae408",
   200 => x"802e81ae",
   201 => x"38bf0baa",
   202 => x"b40cbf0b",
   203 => x"fc0ca8bc",
   204 => x"518dcc2d",
   205 => x"8bb02d87",
   206 => x"f32d8ddc",
   207 => x"2da9a40b",
   208 => x"80f52d70",
   209 => x"872baab4",
   210 => x"08708106",
   211 => x"53565452",
   212 => x"71802e85",
   213 => x"38728107",
   214 => x"5373812a",
   215 => x"70810651",
   216 => x"5271802e",
   217 => x"85387282",
   218 => x"07537382",
   219 => x"2a708106",
   220 => x"51527180",
   221 => x"2e853872",
   222 => x"84075373",
   223 => x"832a7081",
   224 => x"06515271",
   225 => x"802e8538",
   226 => x"72880753",
   227 => x"73842a70",
   228 => x"81065152",
   229 => x"71802e85",
   230 => x"38729007",
   231 => x"5373852a",
   232 => x"70810651",
   233 => x"5271802e",
   234 => x"853872a0",
   235 => x"07537386",
   236 => x"2a708106",
   237 => x"51527180",
   238 => x"2e863872",
   239 => x"80c00753",
   240 => x"72fc0c86",
   241 => x"52aae408",
   242 => x"83388452",
   243 => x"71ec0c86",
   244 => x"b704800b",
   245 => x"aae40c02",
   246 => x"90050d04",
   247 => x"71980c04",
   248 => x"ffb008aa",
   249 => x"e40c0481",
   250 => x"0bffb00c",
   251 => x"04800bff",
   252 => x"b00c0402",
   253 => x"f4050d88",
   254 => x"f504aae4",
   255 => x"0881f02e",
   256 => x"09810689",
   257 => x"38810baa",
   258 => x"ac0c88f5",
   259 => x"04aae408",
   260 => x"81e02e09",
   261 => x"81068938",
   262 => x"810baab0",
   263 => x"0c88f504",
   264 => x"aae40852",
   265 => x"aab00880",
   266 => x"2e8838aa",
   267 => x"e4088180",
   268 => x"05527184",
   269 => x"2c728f06",
   270 => x"5353aaac",
   271 => x"08802e99",
   272 => x"38728429",
   273 => x"a9ec0572",
   274 => x"1381712b",
   275 => x"70097308",
   276 => x"06730c51",
   277 => x"535388eb",
   278 => x"04728429",
   279 => x"a9ec0572",
   280 => x"1383712b",
   281 => x"72080772",
   282 => x"0c535380",
   283 => x"0baab00c",
   284 => x"800baaac",
   285 => x"0cab8051",
   286 => x"89f62daa",
   287 => x"e408ff24",
   288 => x"fef83880",
   289 => x"0baae40c",
   290 => x"028c050d",
   291 => x"0402f805",
   292 => x"0da9ec52",
   293 => x"8f518072",
   294 => x"70840554",
   295 => x"0cff1151",
   296 => x"708025f2",
   297 => x"38028805",
   298 => x"0d0402f0",
   299 => x"050d7551",
   300 => x"87ed2d70",
   301 => x"822cfc06",
   302 => x"a9ec1172",
   303 => x"109e0671",
   304 => x"0870722a",
   305 => x"70830682",
   306 => x"742b7009",
   307 => x"7406760c",
   308 => x"54515657",
   309 => x"53515387",
   310 => x"e72d71aa",
   311 => x"e40c0290",
   312 => x"050d0402",
   313 => x"fc050d72",
   314 => x"5180710c",
   315 => x"800b8412",
   316 => x"0c028405",
   317 => x"0d0402f0",
   318 => x"050d7570",
   319 => x"08841208",
   320 => x"535353ff",
   321 => x"5471712e",
   322 => x"a83887ed",
   323 => x"2d841308",
   324 => x"70842914",
   325 => x"88117008",
   326 => x"7081ff06",
   327 => x"84180881",
   328 => x"11870684",
   329 => x"1a0c5351",
   330 => x"55515151",
   331 => x"87e72d71",
   332 => x"5473aae4",
   333 => x"0c029005",
   334 => x"0d0402f8",
   335 => x"050d87ed",
   336 => x"2de00870",
   337 => x"8b2a7081",
   338 => x"06515252",
   339 => x"70802e9d",
   340 => x"38ab8008",
   341 => x"708429ab",
   342 => x"88057381",
   343 => x"ff06710c",
   344 => x"5151ab80",
   345 => x"08811187",
   346 => x"06ab800c",
   347 => x"51800bab",
   348 => x"a80c87e0",
   349 => x"2d87e72d",
   350 => x"0288050d",
   351 => x"0402fc05",
   352 => x"0d87ed2d",
   353 => x"810baba8",
   354 => x"0c87e72d",
   355 => x"aba80851",
   356 => x"70fa3802",
   357 => x"84050d04",
   358 => x"02fc050d",
   359 => x"ab805189",
   360 => x"e32d898d",
   361 => x"2d8aba51",
   362 => x"87dc2d02",
   363 => x"84050d04",
   364 => x"02fc050d",
   365 => x"810baae0",
   366 => x"0c815184",
   367 => x"8a2d0284",
   368 => x"050d0402",
   369 => x"fc050d8b",
   370 => x"cd0487f3",
   371 => x"2d80f651",
   372 => x"89aa2daa",
   373 => x"e408f338",
   374 => x"80da5189",
   375 => x"aa2daae4",
   376 => x"08e838aa",
   377 => x"dc085189",
   378 => x"aa2daae4",
   379 => x"08dc38aa",
   380 => x"e408aae0",
   381 => x"0caae408",
   382 => x"51848a2d",
   383 => x"0284050d",
   384 => x"0402ec05",
   385 => x"0d765480",
   386 => x"52870b88",
   387 => x"1580f52d",
   388 => x"56537472",
   389 => x"248338a0",
   390 => x"53725182",
   391 => x"f82d8112",
   392 => x"8b1580f5",
   393 => x"2d545272",
   394 => x"7225de38",
   395 => x"0294050d",
   396 => x"0402f005",
   397 => x"0dabb008",
   398 => x"5481f72d",
   399 => x"800babb4",
   400 => x"0c730880",
   401 => x"2e818038",
   402 => x"820baaf8",
   403 => x"0cabb408",
   404 => x"8f06aaf4",
   405 => x"0c730852",
   406 => x"71832e96",
   407 => x"38718326",
   408 => x"89387181",
   409 => x"2eaf388d",
   410 => x"b2047185",
   411 => x"2e9f388d",
   412 => x"b2048814",
   413 => x"80f52d84",
   414 => x"1508a78c",
   415 => x"53545285",
   416 => x"9b2d7184",
   417 => x"29137008",
   418 => x"52528db6",
   419 => x"0473518c",
   420 => x"812d8db2",
   421 => x"04aab408",
   422 => x"8815082c",
   423 => x"70810651",
   424 => x"5271802e",
   425 => x"8738a790",
   426 => x"518daf04",
   427 => x"a7945185",
   428 => x"9b2d8414",
   429 => x"0851859b",
   430 => x"2dabb408",
   431 => x"8105abb4",
   432 => x"0c8c1454",
   433 => x"8cc10402",
   434 => x"90050d04",
   435 => x"71abb00c",
   436 => x"8cb12dab",
   437 => x"b408ff05",
   438 => x"abb80c04",
   439 => x"02e8050d",
   440 => x"abb008ab",
   441 => x"bc085755",
   442 => x"80f65189",
   443 => x"aa2daae4",
   444 => x"08812a70",
   445 => x"81065152",
   446 => x"71802e9f",
   447 => x"388e8304",
   448 => x"87f32d80",
   449 => x"f65189aa",
   450 => x"2daae408",
   451 => x"f338aae0",
   452 => x"08813270",
   453 => x"aae00c51",
   454 => x"848a2d80",
   455 => x"0babac0c",
   456 => x"8c5189aa",
   457 => x"2daae408",
   458 => x"812a7081",
   459 => x"06515271",
   460 => x"802ebf38",
   461 => x"aab808aa",
   462 => x"cc08aab8",
   463 => x"0caacc0c",
   464 => x"aabc08aa",
   465 => x"d008aabc",
   466 => x"0caad00c",
   467 => x"aac008aa",
   468 => x"d408aac0",
   469 => x"0caad40c",
   470 => x"aac408aa",
   471 => x"d808aac4",
   472 => x"0caad80c",
   473 => x"aac808aa",
   474 => x"dc08aac8",
   475 => x"0c70aadc",
   476 => x"0c52aae0",
   477 => x"0881ea38",
   478 => x"aacc0851",
   479 => x"89aa2daa",
   480 => x"e408802e",
   481 => x"8938abac",
   482 => x"088107ab",
   483 => x"ac0caad0",
   484 => x"085189aa",
   485 => x"2daae408",
   486 => x"802e8938",
   487 => x"abac0882",
   488 => x"07abac0c",
   489 => x"aad40851",
   490 => x"89aa2daa",
   491 => x"e408802e",
   492 => x"8938abac",
   493 => x"088407ab",
   494 => x"ac0caad8",
   495 => x"085189aa",
   496 => x"2daae408",
   497 => x"802e8938",
   498 => x"abac0888",
   499 => x"07abac0c",
   500 => x"aadc0851",
   501 => x"89aa2daa",
   502 => x"e408802e",
   503 => x"8938abac",
   504 => x"089007ab",
   505 => x"ac0caab8",
   506 => x"085189aa",
   507 => x"2daae408",
   508 => x"802e8a38",
   509 => x"abac0882",
   510 => x"8007abac",
   511 => x"0caabc08",
   512 => x"5189aa2d",
   513 => x"aae40880",
   514 => x"2e8a38ab",
   515 => x"ac088480",
   516 => x"07abac0c",
   517 => x"aac00851",
   518 => x"89aa2daa",
   519 => x"e408802e",
   520 => x"8a38abac",
   521 => x"08888007",
   522 => x"abac0caa",
   523 => x"c4085189",
   524 => x"aa2daae4",
   525 => x"08802e8a",
   526 => x"38abac08",
   527 => x"908007ab",
   528 => x"ac0caac8",
   529 => x"085189aa",
   530 => x"2daae408",
   531 => x"802e8a38",
   532 => x"abac08a0",
   533 => x"8007abac",
   534 => x"0cabac08",
   535 => x"ed0c96f6",
   536 => x"0481f551",
   537 => x"89aa2daa",
   538 => x"e408812a",
   539 => x"70810651",
   540 => x"52719738",
   541 => x"aacc0851",
   542 => x"89aa2daa",
   543 => x"e408812a",
   544 => x"70810651",
   545 => x"5271802e",
   546 => x"af38abb8",
   547 => x"08527180",
   548 => x"2e8938ff",
   549 => x"12abb80c",
   550 => x"91b804ab",
   551 => x"b40810ab",
   552 => x"b4080570",
   553 => x"84291651",
   554 => x"52881208",
   555 => x"802e8938",
   556 => x"ff518812",
   557 => x"0852712d",
   558 => x"81f25189",
   559 => x"aa2daae4",
   560 => x"08812a70",
   561 => x"81065152",
   562 => x"719738aa",
   563 => x"d0085189",
   564 => x"aa2daae4",
   565 => x"08812a70",
   566 => x"81065152",
   567 => x"71802eb1",
   568 => x"38abb408",
   569 => x"ff11abb8",
   570 => x"08565353",
   571 => x"73722589",
   572 => x"388114ab",
   573 => x"b80c9291",
   574 => x"04721013",
   575 => x"70842916",
   576 => x"51528812",
   577 => x"08802e89",
   578 => x"38fe5188",
   579 => x"12085271",
   580 => x"2d81fd51",
   581 => x"89aa2daa",
   582 => x"e408812a",
   583 => x"70810651",
   584 => x"52719738",
   585 => x"aad40851",
   586 => x"89aa2daa",
   587 => x"e408812a",
   588 => x"70810651",
   589 => x"5271802e",
   590 => x"ad38abb8",
   591 => x"08802e89",
   592 => x"38800bab",
   593 => x"b80c92e6",
   594 => x"04abb408",
   595 => x"10abb408",
   596 => x"05708429",
   597 => x"16515288",
   598 => x"1208802e",
   599 => x"8938fd51",
   600 => x"88120852",
   601 => x"712d81fa",
   602 => x"5189aa2d",
   603 => x"aae40881",
   604 => x"2a708106",
   605 => x"51527197",
   606 => x"38aad808",
   607 => x"5189aa2d",
   608 => x"aae40881",
   609 => x"2a708106",
   610 => x"51527180",
   611 => x"2eae38ab",
   612 => x"b408ff11",
   613 => x"5452abb8",
   614 => x"08732588",
   615 => x"3872abb8",
   616 => x"0c93bc04",
   617 => x"71101270",
   618 => x"84291651",
   619 => x"52881208",
   620 => x"802e8938",
   621 => x"fc518812",
   622 => x"0852712d",
   623 => x"abb80870",
   624 => x"53547380",
   625 => x"2e8a388c",
   626 => x"15ff1555",
   627 => x"5593c204",
   628 => x"820baaf8",
   629 => x"0c718f06",
   630 => x"aaf40c81",
   631 => x"eb5189aa",
   632 => x"2daae408",
   633 => x"812a7081",
   634 => x"06515271",
   635 => x"802ead38",
   636 => x"7408852e",
   637 => x"098106a4",
   638 => x"38881580",
   639 => x"f52dff05",
   640 => x"52718816",
   641 => x"81b72d71",
   642 => x"982b5271",
   643 => x"80258838",
   644 => x"800b8816",
   645 => x"81b72d74",
   646 => x"518c812d",
   647 => x"81f45189",
   648 => x"aa2daae4",
   649 => x"08812a70",
   650 => x"81065152",
   651 => x"71802eb3",
   652 => x"38740885",
   653 => x"2e098106",
   654 => x"aa388815",
   655 => x"80f52d81",
   656 => x"05527188",
   657 => x"1681b72d",
   658 => x"7181ff06",
   659 => x"8b1680f5",
   660 => x"2d545272",
   661 => x"72278738",
   662 => x"72881681",
   663 => x"b72d7451",
   664 => x"8c812d80",
   665 => x"da5189aa",
   666 => x"2daae408",
   667 => x"812a7081",
   668 => x"06515271",
   669 => x"9838aadc",
   670 => x"085189aa",
   671 => x"2daae408",
   672 => x"812a7081",
   673 => x"06515271",
   674 => x"802e81a6",
   675 => x"38abb008",
   676 => x"abb80855",
   677 => x"5373802e",
   678 => x"8a388c13",
   679 => x"ff155553",
   680 => x"95950472",
   681 => x"08527182",
   682 => x"2ea63871",
   683 => x"82268938",
   684 => x"71812ea9",
   685 => x"3896b204",
   686 => x"71832eb1",
   687 => x"3871842e",
   688 => x"09810680",
   689 => x"ed388813",
   690 => x"08518dcc",
   691 => x"2d96b204",
   692 => x"abb80851",
   693 => x"88130852",
   694 => x"712d96b2",
   695 => x"04810b88",
   696 => x"14082baa",
   697 => x"b40832aa",
   698 => x"b40c9688",
   699 => x"04881380",
   700 => x"f52d8105",
   701 => x"8b1480f5",
   702 => x"2d535471",
   703 => x"74248338",
   704 => x"80547388",
   705 => x"1481b72d",
   706 => x"8cb12d96",
   707 => x"b2047508",
   708 => x"802ea238",
   709 => x"75085189",
   710 => x"aa2daae4",
   711 => x"08810652",
   712 => x"71802e8b",
   713 => x"38abb808",
   714 => x"51841608",
   715 => x"52712d88",
   716 => x"165675da",
   717 => x"38805480",
   718 => x"0baaf80c",
   719 => x"738f06aa",
   720 => x"f40ca052",
   721 => x"73abb808",
   722 => x"2e098106",
   723 => x"9838abb4",
   724 => x"08ff0574",
   725 => x"32700981",
   726 => x"05707207",
   727 => x"9f2a9171",
   728 => x"31515153",
   729 => x"53715182",
   730 => x"f82d8114",
   731 => x"548e7425",
   732 => x"c638aae0",
   733 => x"085271aa",
   734 => x"e40c0298",
   735 => x"050d0402",
   736 => x"f4050dd4",
   737 => x"5281ff72",
   738 => x"0c710853",
   739 => x"81ff720c",
   740 => x"72882b83",
   741 => x"fe800672",
   742 => x"087081ff",
   743 => x"06515253",
   744 => x"81ff720c",
   745 => x"72710788",
   746 => x"2b720870",
   747 => x"81ff0651",
   748 => x"525381ff",
   749 => x"720c7271",
   750 => x"07882b72",
   751 => x"087081ff",
   752 => x"067207aa",
   753 => x"e40c5253",
   754 => x"028c050d",
   755 => x"0402f405",
   756 => x"0d747671",
   757 => x"81ff06d4",
   758 => x"0c5353ab",
   759 => x"c0088538",
   760 => x"71892b52",
   761 => x"71982ad4",
   762 => x"0c71902a",
   763 => x"7081ff06",
   764 => x"d40c5171",
   765 => x"882a7081",
   766 => x"ff06d40c",
   767 => x"517181ff",
   768 => x"06d40c72",
   769 => x"902a7081",
   770 => x"ff06d40c",
   771 => x"51d40870",
   772 => x"81ff0651",
   773 => x"5182b8bf",
   774 => x"527081ff",
   775 => x"2e098106",
   776 => x"943881ff",
   777 => x"0bd40cd4",
   778 => x"087081ff",
   779 => x"06ff1454",
   780 => x"515171e5",
   781 => x"3870aae4",
   782 => x"0c028c05",
   783 => x"0d0402fc",
   784 => x"050d81c7",
   785 => x"5181ff0b",
   786 => x"d40cff11",
   787 => x"51708025",
   788 => x"f4380284",
   789 => x"050d0402",
   790 => x"f4050d81",
   791 => x"ff0bd40c",
   792 => x"93538052",
   793 => x"87fc80c1",
   794 => x"5197cd2d",
   795 => x"aae4088b",
   796 => x"3881ff0b",
   797 => x"d40c8153",
   798 => x"99840498",
   799 => x"be2dff13",
   800 => x"5372df38",
   801 => x"72aae40c",
   802 => x"028c050d",
   803 => x"0402ec05",
   804 => x"0d810bab",
   805 => x"c00c8454",
   806 => x"d008708f",
   807 => x"2a708106",
   808 => x"51515372",
   809 => x"f33872d0",
   810 => x"0c98be2d",
   811 => x"a7985185",
   812 => x"9b2dd008",
   813 => x"708f2a70",
   814 => x"81065151",
   815 => x"5372f338",
   816 => x"810bd00c",
   817 => x"b1538052",
   818 => x"84d480c0",
   819 => x"5197cd2d",
   820 => x"aae40881",
   821 => x"2e933872",
   822 => x"822ebd38",
   823 => x"ff135372",
   824 => x"e538ff14",
   825 => x"5473ffb0",
   826 => x"3898be2d",
   827 => x"83aa5284",
   828 => x"9c80c851",
   829 => x"97cd2daa",
   830 => x"e408812e",
   831 => x"09810692",
   832 => x"3896ff2d",
   833 => x"aae40883",
   834 => x"ffff0653",
   835 => x"7283aa2e",
   836 => x"9d3898d7",
   837 => x"2d9aa904",
   838 => x"a7a45185",
   839 => x"9b2d8053",
   840 => x"9bf704a7",
   841 => x"bc51859b",
   842 => x"2d80549b",
   843 => x"c90481ff",
   844 => x"0bd40cb1",
   845 => x"5498be2d",
   846 => x"8fcf5380",
   847 => x"5287fc80",
   848 => x"f75197cd",
   849 => x"2daae408",
   850 => x"55aae408",
   851 => x"812e0981",
   852 => x"069b3881",
   853 => x"ff0bd40c",
   854 => x"820a5284",
   855 => x"9c80e951",
   856 => x"97cd2daa",
   857 => x"e408802e",
   858 => x"8d3898be",
   859 => x"2dff1353",
   860 => x"72c9389b",
   861 => x"bc0481ff",
   862 => x"0bd40caa",
   863 => x"e4085287",
   864 => x"fc80fa51",
   865 => x"97cd2daa",
   866 => x"e408b138",
   867 => x"81ff0bd4",
   868 => x"0cd40853",
   869 => x"81ff0bd4",
   870 => x"0c81ff0b",
   871 => x"d40c81ff",
   872 => x"0bd40c81",
   873 => x"ff0bd40c",
   874 => x"72862a70",
   875 => x"81067656",
   876 => x"51537295",
   877 => x"38aae408",
   878 => x"549bc904",
   879 => x"73822efe",
   880 => x"e238ff14",
   881 => x"5473feed",
   882 => x"3873abc0",
   883 => x"0c738b38",
   884 => x"815287fc",
   885 => x"80d05197",
   886 => x"cd2d81ff",
   887 => x"0bd40cd0",
   888 => x"08708f2a",
   889 => x"70810651",
   890 => x"515372f3",
   891 => x"3872d00c",
   892 => x"81ff0bd4",
   893 => x"0c815372",
   894 => x"aae40c02",
   895 => x"94050d04",
   896 => x"02e8050d",
   897 => x"78558056",
   898 => x"81ff0bd4",
   899 => x"0cd00870",
   900 => x"8f2a7081",
   901 => x"06515153",
   902 => x"72f33882",
   903 => x"810bd00c",
   904 => x"81ff0bd4",
   905 => x"0c775287",
   906 => x"fc80d151",
   907 => x"97cd2d80",
   908 => x"dbc6df54",
   909 => x"aae40880",
   910 => x"2e8a38a7",
   911 => x"dc51859b",
   912 => x"2d9d9704",
   913 => x"81ff0bd4",
   914 => x"0cd40870",
   915 => x"81ff0651",
   916 => x"537281fe",
   917 => x"2e098106",
   918 => x"9d3880ff",
   919 => x"5396ff2d",
   920 => x"aae40875",
   921 => x"70840557",
   922 => x"0cff1353",
   923 => x"728025ed",
   924 => x"3881569c",
   925 => x"fc04ff14",
   926 => x"5473c938",
   927 => x"81ff0bd4",
   928 => x"0c81ff0b",
   929 => x"d40cd008",
   930 => x"708f2a70",
   931 => x"81065151",
   932 => x"5372f338",
   933 => x"72d00c75",
   934 => x"aae40c02",
   935 => x"98050d04",
   936 => x"02e8050d",
   937 => x"77797b58",
   938 => x"55558053",
   939 => x"727625a3",
   940 => x"38747081",
   941 => x"055680f5",
   942 => x"2d747081",
   943 => x"055680f5",
   944 => x"2d525271",
   945 => x"712e8638",
   946 => x"81519dd5",
   947 => x"04811353",
   948 => x"9dac0480",
   949 => x"5170aae4",
   950 => x"0c029805",
   951 => x"0d0402ec",
   952 => x"050d7655",
   953 => x"74802ebb",
   954 => x"389a1580",
   955 => x"e02d51a4",
   956 => x"e22daae4",
   957 => x"08aae408",
   958 => x"aff00caa",
   959 => x"e4085454",
   960 => x"afcc0880",
   961 => x"2e993894",
   962 => x"1580e02d",
   963 => x"51a4e22d",
   964 => x"aae40890",
   965 => x"2b83fff0",
   966 => x"0a067075",
   967 => x"07515372",
   968 => x"aff00caf",
   969 => x"f0085372",
   970 => x"802e9938",
   971 => x"afc408fe",
   972 => x"147129af",
   973 => x"d80805af",
   974 => x"f40c7084",
   975 => x"2bafd00c",
   976 => x"549eea04",
   977 => x"afdc08af",
   978 => x"f00cafe0",
   979 => x"08aff40c",
   980 => x"afcc0880",
   981 => x"2e8a38af",
   982 => x"c408842b",
   983 => x"539ee604",
   984 => x"afe40884",
   985 => x"2b5372af",
   986 => x"d00c0294",
   987 => x"050d0402",
   988 => x"d8050d80",
   989 => x"0bafcc0c",
   990 => x"8454998d",
   991 => x"2daae408",
   992 => x"802e9538",
   993 => x"abc45280",
   994 => x"519c802d",
   995 => x"aae40880",
   996 => x"2e8638fe",
   997 => x"549fa004",
   998 => x"ff145473",
   999 => x"8024db38",
  1000 => x"738c38a7",
  1001 => x"ec51859b",
  1002 => x"2d7355a4",
  1003 => x"a9048056",
  1004 => x"810baff8",
  1005 => x"0c8853a8",
  1006 => x"8052abfa",
  1007 => x"519da02d",
  1008 => x"aae40876",
  1009 => x"2e098106",
  1010 => x"8738aae4",
  1011 => x"08aff80c",
  1012 => x"8853a88c",
  1013 => x"52ac9651",
  1014 => x"9da02daa",
  1015 => x"e4088738",
  1016 => x"aae408af",
  1017 => x"f80caff8",
  1018 => x"08802e80",
  1019 => x"f638af8a",
  1020 => x"0b80f52d",
  1021 => x"af8b0b80",
  1022 => x"f52d7198",
  1023 => x"2b71902b",
  1024 => x"07af8c0b",
  1025 => x"80f52d70",
  1026 => x"882b7207",
  1027 => x"af8d0b80",
  1028 => x"f52d7107",
  1029 => x"afc20b80",
  1030 => x"f52dafc3",
  1031 => x"0b80f52d",
  1032 => x"71882b07",
  1033 => x"535f5452",
  1034 => x"5a565755",
  1035 => x"7381abaa",
  1036 => x"2e098106",
  1037 => x"8d387551",
  1038 => x"a4b22daa",
  1039 => x"e40856a0",
  1040 => x"cf047382",
  1041 => x"d4d52e87",
  1042 => x"38a89851",
  1043 => x"a19004ab",
  1044 => x"c4527551",
  1045 => x"9c802daa",
  1046 => x"e40855aa",
  1047 => x"e408802e",
  1048 => x"83c73888",
  1049 => x"53a88c52",
  1050 => x"ac96519d",
  1051 => x"a02daae4",
  1052 => x"08893881",
  1053 => x"0bafcc0c",
  1054 => x"a1960488",
  1055 => x"53a88052",
  1056 => x"abfa519d",
  1057 => x"a02daae4",
  1058 => x"08802e8a",
  1059 => x"38a8ac51",
  1060 => x"859b2da1",
  1061 => x"f004afc2",
  1062 => x"0b80f52d",
  1063 => x"547380d5",
  1064 => x"2e098106",
  1065 => x"80ca38af",
  1066 => x"c30b80f5",
  1067 => x"2d547381",
  1068 => x"aa2e0981",
  1069 => x"06ba3880",
  1070 => x"0babc40b",
  1071 => x"80f52d56",
  1072 => x"547481e9",
  1073 => x"2e833881",
  1074 => x"547481eb",
  1075 => x"2e8c3880",
  1076 => x"5573752e",
  1077 => x"09810682",
  1078 => x"d038abcf",
  1079 => x"0b80f52d",
  1080 => x"55748d38",
  1081 => x"abd00b80",
  1082 => x"f52d5473",
  1083 => x"822e8638",
  1084 => x"8055a4a9",
  1085 => x"04abd10b",
  1086 => x"80f52d70",
  1087 => x"afc40cff",
  1088 => x"05afc80c",
  1089 => x"abd20b80",
  1090 => x"f52dabd3",
  1091 => x"0b80f52d",
  1092 => x"58760577",
  1093 => x"82802905",
  1094 => x"70afd40c",
  1095 => x"abd40b80",
  1096 => x"f52d70af",
  1097 => x"e80cafcc",
  1098 => x"08595758",
  1099 => x"76802e81",
  1100 => x"a3388853",
  1101 => x"a88c52ac",
  1102 => x"96519da0",
  1103 => x"2daae408",
  1104 => x"81e738af",
  1105 => x"c4087084",
  1106 => x"2bafd00c",
  1107 => x"70afe40c",
  1108 => x"abe90b80",
  1109 => x"f52dabe8",
  1110 => x"0b80f52d",
  1111 => x"71828029",
  1112 => x"05abea0b",
  1113 => x"80f52d70",
  1114 => x"84808029",
  1115 => x"12abeb0b",
  1116 => x"80f52d70",
  1117 => x"81800a29",
  1118 => x"1270afec",
  1119 => x"0cafe808",
  1120 => x"7129afd4",
  1121 => x"080570af",
  1122 => x"d80cabf1",
  1123 => x"0b80f52d",
  1124 => x"abf00b80",
  1125 => x"f52d7182",
  1126 => x"802905ab",
  1127 => x"f20b80f5",
  1128 => x"2d708480",
  1129 => x"802912ab",
  1130 => x"f30b80f5",
  1131 => x"2d70982b",
  1132 => x"81f00a06",
  1133 => x"720570af",
  1134 => x"dc0cfe11",
  1135 => x"7e297705",
  1136 => x"afe00c52",
  1137 => x"59524354",
  1138 => x"5e515259",
  1139 => x"525d5759",
  1140 => x"57a4a204",
  1141 => x"abd60b80",
  1142 => x"f52dabd5",
  1143 => x"0b80f52d",
  1144 => x"71828029",
  1145 => x"0570afd0",
  1146 => x"0c70a029",
  1147 => x"83ff0570",
  1148 => x"892a70af",
  1149 => x"e40cabdb",
  1150 => x"0b80f52d",
  1151 => x"abda0b80",
  1152 => x"f52d7182",
  1153 => x"80290570",
  1154 => x"afec0c7b",
  1155 => x"71291e70",
  1156 => x"afe00c7d",
  1157 => x"afdc0c73",
  1158 => x"05afd80c",
  1159 => x"555e5151",
  1160 => x"55558051",
  1161 => x"9dde2d81",
  1162 => x"5574aae4",
  1163 => x"0c02a805",
  1164 => x"0d0402f4",
  1165 => x"050d7470",
  1166 => x"882a83fe",
  1167 => x"80067072",
  1168 => x"982a0772",
  1169 => x"882b87fc",
  1170 => x"80800673",
  1171 => x"982b81f0",
  1172 => x"0a067173",
  1173 => x"0707aae4",
  1174 => x"0c565153",
  1175 => x"51028c05",
  1176 => x"0d0402f8",
  1177 => x"050d028e",
  1178 => x"0580f52d",
  1179 => x"74882b07",
  1180 => x"7083ffff",
  1181 => x"06aae40c",
  1182 => x"51028805",
  1183 => x"0d040000",
  1184 => x"00ffffff",
  1185 => x"ff00ffff",
  1186 => x"ffff00ff",
  1187 => x"ffffff00",
  1188 => x"52657365",
  1189 => x"74000000",
  1190 => x"4d616e75",
  1191 => x"616c2053",
  1192 => x"65727665",
  1193 => x"00000000",
  1194 => x"42616c6c",
  1195 => x"20416e67",
  1196 => x"6c650000",
  1197 => x"42616c6c",
  1198 => x"20537065",
  1199 => x"65640000",
  1200 => x"50616464",
  1201 => x"6c652053",
  1202 => x"697a6500",
  1203 => x"536f756e",
  1204 => x"64000000",
  1205 => x"466f7572",
  1206 => x"20706c61",
  1207 => x"79657273",
  1208 => x"00000000",
  1209 => x"446f7562",
  1210 => x"6c65204f",
  1211 => x"53442077",
  1212 => x"696e646f",
  1213 => x"77000000",
  1214 => x"45786974",
  1215 => x"00000000",
  1216 => x"4d6f6e6f",
  1217 => x"00000000",
  1218 => x"47726579",
  1219 => x"7363616c",
  1220 => x"65000000",
  1221 => x"52474231",
  1222 => x"00000000",
  1223 => x"52474232",
  1224 => x"00000000",
  1225 => x"4669656c",
  1226 => x"64000000",
  1227 => x"49636500",
  1228 => x"43687269",
  1229 => x"73746d61",
  1230 => x"73000000",
  1231 => x"4d61726b",
  1232 => x"736d616e",
  1233 => x"00000000",
  1234 => x"4c617320",
  1235 => x"56656761",
  1236 => x"73000000",
  1237 => x"41592d33",
  1238 => x"2d383531",
  1239 => x"3520636f",
  1240 => x"6c6f7273",
  1241 => x"00000000",
  1242 => x"54525120",
  1243 => x"436f6c6f",
  1244 => x"72730000",
  1245 => x"496e6974",
  1246 => x"69616c69",
  1247 => x"7a696e67",
  1248 => x"20534420",
  1249 => x"63617264",
  1250 => x"0a000000",
  1251 => x"16200000",
  1252 => x"14200000",
  1253 => x"15200000",
  1254 => x"53442069",
  1255 => x"6e69742e",
  1256 => x"2e2e0a00",
  1257 => x"53442063",
  1258 => x"61726420",
  1259 => x"72657365",
  1260 => x"74206661",
  1261 => x"696c6564",
  1262 => x"210a0000",
  1263 => x"53444843",
  1264 => x"20657272",
  1265 => x"6f72210a",
  1266 => x"00000000",
  1267 => x"57726974",
  1268 => x"65206661",
  1269 => x"696c6564",
  1270 => x"0a000000",
  1271 => x"52656164",
  1272 => x"20666169",
  1273 => x"6c65640a",
  1274 => x"00000000",
  1275 => x"43617264",
  1276 => x"20696e69",
  1277 => x"74206661",
  1278 => x"696c6564",
  1279 => x"0a000000",
  1280 => x"46415431",
  1281 => x"36202020",
  1282 => x"00000000",
  1283 => x"46415433",
  1284 => x"32202020",
  1285 => x"00000000",
  1286 => x"4e6f2070",
  1287 => x"61727469",
  1288 => x"74696f6e",
  1289 => x"20736967",
  1290 => x"0a000000",
  1291 => x"42616420",
  1292 => x"70617274",
  1293 => x"0a000000",
  1294 => x"00000002",
  1295 => x"00000002",
  1296 => x"00001290",
  1297 => x"000002d4",
  1298 => x"00000001",
  1299 => x"00001298",
  1300 => x"00000000",
  1301 => x"00000001",
  1302 => x"000012a8",
  1303 => x"00000001",
  1304 => x"00000001",
  1305 => x"000012b4",
  1306 => x"00000002",
  1307 => x"00000001",
  1308 => x"000012c0",
  1309 => x"00000003",
  1310 => x"00000001",
  1311 => x"000012cc",
  1312 => x"00000004",
  1313 => x"00000001",
  1314 => x"000012d4",
  1315 => x"00000006",
  1316 => x"00000001",
  1317 => x"000012e4",
  1318 => x"00000005",
  1319 => x"00000003",
  1320 => x"000014c0",
  1321 => x"0000000b",
  1322 => x"00000002",
  1323 => x"000012f8",
  1324 => x"000005c3",
  1325 => x"00000000",
  1326 => x"00000000",
  1327 => x"00000000",
  1328 => x"00001300",
  1329 => x"00001308",
  1330 => x"00001314",
  1331 => x"0000131c",
  1332 => x"00001324",
  1333 => x"0000132c",
  1334 => x"00001330",
  1335 => x"0000133c",
  1336 => x"00001348",
  1337 => x"00001354",
  1338 => x"00001368",
  1339 => x"00000000",
  1340 => x"00000000",
  1341 => x"00000000",
  1342 => x"00000000",
  1343 => x"00000000",
  1344 => x"00000000",
  1345 => x"00000000",
  1346 => x"00000000",
  1347 => x"00000000",
  1348 => x"00000000",
  1349 => x"00000000",
  1350 => x"00000000",
  1351 => x"00000000",
  1352 => x"00000000",
  1353 => x"00000000",
  1354 => x"00000000",
  1355 => x"00000000",
  1356 => x"00000000",
  1357 => x"00000006",
  1358 => x"00000043",
  1359 => x"00000042",
  1360 => x"0000003b",
  1361 => x"0000004b",
  1362 => x"00000033",
  1363 => x"00000003",
  1364 => x"0000000b",
  1365 => x"00000083",
  1366 => x"00000023",
  1367 => x"0000002b",
  1368 => x"00000000",
	others => x"00000000"
);

begin

process (clk)
begin
	if (clk'event and clk = '1') then
		if (from_zpu.memAWriteEnable = '1') and (from_zpu.memBWriteEnable = '1') and (from_zpu.memAAddr=from_zpu.memBAddr) and (from_zpu.memAWrite/=from_zpu.memBWrite) then
			report "write collision" severity failure;
		end if;
	
		if (from_zpu.memAWriteEnable = '1') then
			ram(to_integer(unsigned(from_zpu.memAAddr(maxAddrBitBRAM downto 2)))) := from_zpu.memAWrite;
			to_zpu.memARead <= from_zpu.memAWrite;
		else
			to_zpu.memARead <= ram(to_integer(unsigned(from_zpu.memAAddr(maxAddrBitBRAM downto 2))));
		end if;
	end if;
end process;

process (clk)
begin
	if (clk'event and clk = '1') then
		if (from_zpu.memBWriteEnable = '1') then
			ram(to_integer(unsigned(from_zpu.memBAddr(maxAddrBitBRAM downto 2)))) := from_zpu.memBWrite;
			to_zpu.memBRead <= from_zpu.memBWrite;
		else
			to_zpu.memBRead <= ram(to_integer(unsigned(from_zpu.memBAddr(maxAddrBitBRAM downto 2))));
		end if;
	end if;
end process;


end arch;

