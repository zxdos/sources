library IEEE;
use IEEE.std_logic_1164.all;
use IEEE.numeric_std.all;

entity ROM81hh is
	port(
		Clk	: in std_logic;
		AIn	: in std_logic_vector(11 downto 0);
		D	: out std_logic_vector(7 downto 0)
	);
end ROM81hh;

architecture rtl of ROM81hh is
	signal A	: std_logic_vector(12 downto 0);
begin
	A(10 downto 0) <= AIn(10 downto 0);
	A(12 downto 11) <= "11";
	process (A)
	begin
		case to_integer(unsigned(A)) is
		when 006144 => D <= "00011111";	-- 0x1800
		when 006145 => D <= "00010000";	-- 0x1801
		when 006146 => D <= "11100100";	-- 0x1802
		when 006147 => D <= "11101011";	-- 0x1803
		when 006148 => D <= "11011001";	-- 0x1804
		when 006149 => D <= "11101011";	-- 0x1805
		when 006150 => D <= "11011001";	-- 0x1806
		when 006151 => D <= "11000001";	-- 0x1807
		when 006152 => D <= "11100001";	-- 0x1808
		when 006153 => D <= "01111000";	-- 0x1809
		when 006154 => D <= "10000001";	-- 0x180A
		when 006155 => D <= "00100000";	-- 0x180B
		when 006156 => D <= "00000001";	-- 0x180C
		when 006157 => D <= "10100111";	-- 0x180D
		when 006158 => D <= "00111101";	-- 0x180E
		when 006159 => D <= "00111111";	-- 0x180F
		when 006160 => D <= "00010111";	-- 0x1810
		when 006161 => D <= "00111111";	-- 0x1811
		when 006162 => D <= "00011111";	-- 0x1812
		when 006163 => D <= "11110010";	-- 0x1813
		when 006164 => D <= "00011001";	-- 0x1814
		when 006165 => D <= "00011000";	-- 0x1815
		when 006166 => D <= "00110000";	-- 0x1816
		when 006167 => D <= "01101000";	-- 0x1817
		when 006168 => D <= "10100111";	-- 0x1818
		when 006169 => D <= "00111100";	-- 0x1819
		when 006170 => D <= "00100000";	-- 0x181A
		when 006171 => D <= "00001000";	-- 0x181B
		when 006172 => D <= "00111000";	-- 0x181C
		when 006173 => D <= "00000110";	-- 0x181D
		when 006174 => D <= "11011001";	-- 0x181E
		when 006175 => D <= "11001011";	-- 0x181F
		when 006176 => D <= "01111010";	-- 0x1820
		when 006177 => D <= "11011001";	-- 0x1821
		when 006178 => D <= "00100000";	-- 0x1822
		when 006179 => D <= "01011100";	-- 0x1823
		when 006180 => D <= "01110111";	-- 0x1824
		when 006181 => D <= "11011001";	-- 0x1825
		when 006182 => D <= "01111000";	-- 0x1826
		when 006183 => D <= "11011001";	-- 0x1827
		when 006184 => D <= "00110000";	-- 0x1828
		when 006185 => D <= "00010101";	-- 0x1829
		when 006186 => D <= "01111110";	-- 0x182A
		when 006187 => D <= "10100111";	-- 0x182B
		when 006188 => D <= "00111110";	-- 0x182C
		when 006189 => D <= "10000000";	-- 0x182D
		when 006190 => D <= "00101000";	-- 0x182E
		when 006191 => D <= "00000001";	-- 0x182F
		when 006192 => D <= "10101111";	-- 0x1830
		when 006193 => D <= "11011001";	-- 0x1831
		when 006194 => D <= "10100010";	-- 0x1832
		when 006195 => D <= "11001101";	-- 0x1833
		when 006196 => D <= "00111000";	-- 0x1834
		when 006197 => D <= "00010111";	-- 0x1835
		when 006198 => D <= "00000111";	-- 0x1836
		when 006199 => D <= "01110111";	-- 0x1837
		when 006200 => D <= "00111000";	-- 0x1838
		when 006201 => D <= "00101110";	-- 0x1839
		when 006202 => D <= "00100011";	-- 0x183A
		when 006203 => D <= "01110111";	-- 0x183B
		when 006204 => D <= "00101011";	-- 0x183C
		when 006205 => D <= "00011000";	-- 0x183D
		when 006206 => D <= "00101001";	-- 0x183E
		when 006207 => D <= "00000110";	-- 0x183F
		when 006208 => D <= "00100000";	-- 0x1840
		when 006209 => D <= "11011001";	-- 0x1841
		when 006210 => D <= "11001011";	-- 0x1842
		when 006211 => D <= "01111010";	-- 0x1843
		when 006212 => D <= "11011001";	-- 0x1844
		when 006213 => D <= "00100000";	-- 0x1845
		when 006214 => D <= "00010010";	-- 0x1846
		when 006215 => D <= "00000111";	-- 0x1847
		when 006216 => D <= "11001011";	-- 0x1848
		when 006217 => D <= "00010011";	-- 0x1849
		when 006218 => D <= "11001011";	-- 0x184A
		when 006219 => D <= "00010010";	-- 0x184B
		when 006220 => D <= "11011001";	-- 0x184C
		when 006221 => D <= "11001011";	-- 0x184D
		when 006222 => D <= "00010011";	-- 0x184E
		when 006223 => D <= "11001011";	-- 0x184F
		when 006224 => D <= "00010010";	-- 0x1850
		when 006225 => D <= "11011001";	-- 0x1851
		when 006226 => D <= "00110101";	-- 0x1852
		when 006227 => D <= "00101000";	-- 0x1853
		when 006228 => D <= "11010111";	-- 0x1854
		when 006229 => D <= "00010000";	-- 0x1855
		when 006230 => D <= "11101010";	-- 0x1856
		when 006231 => D <= "00011000";	-- 0x1857
		when 006232 => D <= "11010111";	-- 0x1858
		when 006233 => D <= "00010111";	-- 0x1859
		when 006234 => D <= "00110000";	-- 0x185A
		when 006235 => D <= "00001100";	-- 0x185B
		when 006236 => D <= "11001101";	-- 0x185C
		when 006237 => D <= "01000001";	-- 0x185D
		when 006238 => D <= "00010111";	-- 0x185E
		when 006239 => D <= "00100000";	-- 0x185F
		when 006240 => D <= "00000111";	-- 0x1860
		when 006241 => D <= "11011001";	-- 0x1861
		when 006242 => D <= "00010110";	-- 0x1862
		when 006243 => D <= "10000000";	-- 0x1863
		when 006244 => D <= "11011001";	-- 0x1864
		when 006245 => D <= "00110100";	-- 0x1865
		when 006246 => D <= "00101000";	-- 0x1866
		when 006247 => D <= "00011000";	-- 0x1867
		when 006248 => D <= "11100101";	-- 0x1868
		when 006249 => D <= "00100011";	-- 0x1869
		when 006250 => D <= "11011001";	-- 0x186A
		when 006251 => D <= "11010101";	-- 0x186B
		when 006252 => D <= "11011001";	-- 0x186C
		when 006253 => D <= "11000001";	-- 0x186D
		when 006254 => D <= "01111000";	-- 0x186E
		when 006255 => D <= "00010111";	-- 0x186F
		when 006256 => D <= "11001011";	-- 0x1870
		when 006257 => D <= "00010110";	-- 0x1871
		when 006258 => D <= "00011111";	-- 0x1872
		when 006259 => D <= "01110111";	-- 0x1873
		when 006260 => D <= "00100011";	-- 0x1874
		when 006261 => D <= "01110001";	-- 0x1875
		when 006262 => D <= "00100011";	-- 0x1876
		when 006263 => D <= "01110010";	-- 0x1877
		when 006264 => D <= "00100011";	-- 0x1878
		when 006265 => D <= "01110011";	-- 0x1879
		when 006266 => D <= "11100001";	-- 0x187A
		when 006267 => D <= "11010001";	-- 0x187B
		when 006268 => D <= "11011001";	-- 0x187C
		when 006269 => D <= "11100001";	-- 0x187D
		when 006270 => D <= "11011001";	-- 0x187E
		when 006271 => D <= "11001001";	-- 0x187F
		when 006272 => D <= "11001111";	-- 0x1880
		when 006273 => D <= "00000101";	-- 0x1881
		when 006274 => D <= "11101011";	-- 0x1882
		when 006275 => D <= "10101111";	-- 0x1883
		when 006276 => D <= "11001101";	-- 0x1884
		when 006277 => D <= "10111100";	-- 0x1885
		when 006278 => D <= "00010111";	-- 0x1886
		when 006279 => D <= "00111000";	-- 0x1887
		when 006280 => D <= "11110111";	-- 0x1888
		when 006281 => D <= "11101011";	-- 0x1889
		when 006282 => D <= "11001101";	-- 0x188A
		when 006283 => D <= "10111100";	-- 0x188B
		when 006284 => D <= "00010111";	-- 0x188C
		when 006285 => D <= "11011000";	-- 0x188D
		when 006286 => D <= "11011001";	-- 0x188E
		when 006287 => D <= "11100101";	-- 0x188F
		when 006288 => D <= "11011001";	-- 0x1890
		when 006289 => D <= "11010101";	-- 0x1891
		when 006290 => D <= "11100101";	-- 0x1892
		when 006291 => D <= "11001101";	-- 0x1893
		when 006292 => D <= "11110111";	-- 0x1894
		when 006293 => D <= "00010110";	-- 0x1895
		when 006294 => D <= "11011001";	-- 0x1896
		when 006295 => D <= "11100101";	-- 0x1897
		when 006296 => D <= "01100000";	-- 0x1898
		when 006297 => D <= "01101001";	-- 0x1899
		when 006298 => D <= "11011001";	-- 0x189A
		when 006299 => D <= "01100001";	-- 0x189B
		when 006300 => D <= "01101000";	-- 0x189C
		when 006301 => D <= "10101111";	-- 0x189D
		when 006302 => D <= "00000110";	-- 0x189E
		when 006303 => D <= "11011111";	-- 0x189F
		when 006304 => D <= "00011000";	-- 0x18A0
		when 006305 => D <= "00010000";	-- 0x18A1
		when 006306 => D <= "00010111";	-- 0x18A2
		when 006307 => D <= "11001011";	-- 0x18A3
		when 006308 => D <= "00010001";	-- 0x18A4
		when 006309 => D <= "11011001";	-- 0x18A5
		when 006310 => D <= "11001011";	-- 0x18A6
		when 006311 => D <= "00010001";	-- 0x18A7
		when 006312 => D <= "11001011";	-- 0x18A8
		when 006313 => D <= "00010000";	-- 0x18A9
		when 006314 => D <= "11011001";	-- 0x18AA
		when 006315 => D <= "00101001";	-- 0x18AB
		when 006316 => D <= "11011001";	-- 0x18AC
		when 006317 => D <= "11101101";	-- 0x18AD
		when 006318 => D <= "01101010";	-- 0x18AE
		when 006319 => D <= "11011001";	-- 0x18AF
		when 006320 => D <= "00111000";	-- 0x18B0
		when 006321 => D <= "00010000";	-- 0x18B1
		when 006322 => D <= "11101101";	-- 0x18B2
		when 006323 => D <= "01010010";	-- 0x18B3
		when 006324 => D <= "11011001";	-- 0x18B4
		when 006325 => D <= "11101101";	-- 0x18B5
		when 006326 => D <= "01010010";	-- 0x18B6
		when 006327 => D <= "11011001";	-- 0x18B7
		when 006328 => D <= "00110000";	-- 0x18B8
		when 006329 => D <= "00001111";	-- 0x18B9
		when 006330 => D <= "00011001";	-- 0x18BA
		when 006331 => D <= "11011001";	-- 0x18BB
		when 006332 => D <= "11101101";	-- 0x18BC
		when 006333 => D <= "01011010";	-- 0x18BD
		when 006334 => D <= "11011001";	-- 0x18BE
		when 006335 => D <= "10100111";	-- 0x18BF
		when 006336 => D <= "00011000";	-- 0x18C0
		when 006337 => D <= "00001000";	-- 0x18C1
		when 006338 => D <= "10100111";	-- 0x18C2
		when 006339 => D <= "11101101";	-- 0x18C3
		when 006340 => D <= "01010010";	-- 0x18C4
		when 006341 => D <= "11011001";	-- 0x18C5
		when 006342 => D <= "11101101";	-- 0x18C6
		when 006343 => D <= "01010010";	-- 0x18C7
		when 006344 => D <= "11011001";	-- 0x18C8
		when 006345 => D <= "00110111";	-- 0x18C9
		when 006346 => D <= "00000100";	-- 0x18CA
		when 006347 => D <= "11111010";	-- 0x18CB
		when 006348 => D <= "10100010";	-- 0x18CC
		when 006349 => D <= "00011000";	-- 0x18CD
		when 006350 => D <= "11110101";	-- 0x18CE
		when 006351 => D <= "00101000";	-- 0x18CF
		when 006352 => D <= "11100001";	-- 0x18D0
		when 006353 => D <= "01011111";	-- 0x18D1
		when 006354 => D <= "01010001";	-- 0x18D2
		when 006355 => D <= "11011001";	-- 0x18D3
		when 006356 => D <= "01011001";	-- 0x18D4
		when 006357 => D <= "01010000";	-- 0x18D5
		when 006358 => D <= "11110001";	-- 0x18D6
		when 006359 => D <= "11001011";	-- 0x18D7
		when 006360 => D <= "00011000";	-- 0x18D8
		when 006361 => D <= "11110001";	-- 0x18D9
		when 006362 => D <= "11001011";	-- 0x18DA
		when 006363 => D <= "00011000";	-- 0x18DB
		when 006364 => D <= "11011001";	-- 0x18DC
		when 006365 => D <= "11000001";	-- 0x18DD
		when 006366 => D <= "11100001";	-- 0x18DE
		when 006367 => D <= "01111000";	-- 0x18DF
		when 006368 => D <= "10010001";	-- 0x18E0
		when 006369 => D <= "11000011";	-- 0x18E1
		when 006370 => D <= "00010000";	-- 0x18E2
		when 006371 => D <= "00011000";	-- 0x18E3
		when 006372 => D <= "01111110";	-- 0x18E4
		when 006373 => D <= "11111110";	-- 0x18E5
		when 006374 => D <= "10000001";	-- 0x18E6
		when 006375 => D <= "00110000";	-- 0x18E7
		when 006376 => D <= "00000110";	-- 0x18E8
		when 006377 => D <= "00110110";	-- 0x18E9
		when 006378 => D <= "00000000";	-- 0x18EA
		when 006379 => D <= "00111110";	-- 0x18EB
		when 006380 => D <= "00100000";	-- 0x18EC
		when 006381 => D <= "00011000";	-- 0x18ED
		when 006382 => D <= "00000101";	-- 0x18EE
		when 006383 => D <= "11010110";	-- 0x18EF
		when 006384 => D <= "10100000";	-- 0x18F0
		when 006385 => D <= "11110000";	-- 0x18F1
		when 006386 => D <= "11101101";	-- 0x18F2
		when 006387 => D <= "01000100";	-- 0x18F3
		when 006388 => D <= "11010101";	-- 0x18F4
		when 006389 => D <= "11101011";	-- 0x18F5
		when 006390 => D <= "00101011";	-- 0x18F6
		when 006391 => D <= "01000111";	-- 0x18F7
		when 006392 => D <= "11001011";	-- 0x18F8
		when 006393 => D <= "00111000";	-- 0x18F9
		when 006394 => D <= "11001011";	-- 0x18FA
		when 006395 => D <= "00111000";	-- 0x18FB
		when 006396 => D <= "11001011";	-- 0x18FC
		when 006397 => D <= "00111000";	-- 0x18FD
		when 006398 => D <= "00101000";	-- 0x18FE
		when 006399 => D <= "00000101";	-- 0x18FF
		when 006400 => D <= "00110110";	-- 0x1900
		when 006401 => D <= "00000000";	-- 0x1901
		when 006402 => D <= "00101011";	-- 0x1902
		when 006403 => D <= "00010000";	-- 0x1903
		when 006404 => D <= "11111011";	-- 0x1904
		when 006405 => D <= "11100110";	-- 0x1905
		when 006406 => D <= "00000111";	-- 0x1906
		when 006407 => D <= "00101000";	-- 0x1907
		when 006408 => D <= "00001001";	-- 0x1908
		when 006409 => D <= "01000111";	-- 0x1909
		when 006410 => D <= "00111110";	-- 0x190A
		when 006411 => D <= "11111111";	-- 0x190B
		when 006412 => D <= "11001011";	-- 0x190C
		when 006413 => D <= "00100111";	-- 0x190D
		when 006414 => D <= "00010000";	-- 0x190E
		when 006415 => D <= "11111100";	-- 0x190F
		when 006416 => D <= "10100110";	-- 0x1910
		when 006417 => D <= "01110111";	-- 0x1911
		when 006418 => D <= "11101011";	-- 0x1912
		when 006419 => D <= "11010001";	-- 0x1913
		when 006420 => D <= "11001001";	-- 0x1914
		when 006421 => D <= "00000000";	-- 0x1915
		when 006422 => D <= "10110000";	-- 0x1916
		when 006423 => D <= "00000000";	-- 0x1917
		when 006424 => D <= "00110001";	-- 0x1918
		when 006425 => D <= "00000000";	-- 0x1919
		when 006426 => D <= "00110000";	-- 0x191A
		when 006427 => D <= "00000000";	-- 0x191B
		when 006428 => D <= "11110001";	-- 0x191C
		when 006429 => D <= "01001001";	-- 0x191D
		when 006430 => D <= "00001111";	-- 0x191E
		when 006431 => D <= "11011010";	-- 0x191F
		when 006432 => D <= "10100010";	-- 0x1920
		when 006433 => D <= "00110100";	-- 0x1921
		when 006434 => D <= "00100000";	-- 0x1922
		when 006435 => D <= "00101111";	-- 0x1923
		when 006436 => D <= "00011100";	-- 0x1924
		when 006437 => D <= "01110010";	-- 0x1925
		when 006438 => D <= "00011010";	-- 0x1926
		when 006439 => D <= "11100011";	-- 0x1927
		when 006440 => D <= "00011001";	-- 0x1928
		when 006441 => D <= "01001100";	-- 0x1929
		when 006442 => D <= "00010111";	-- 0x192A
		when 006443 => D <= "11000110";	-- 0x192B
		when 006444 => D <= "00010111";	-- 0x192C
		when 006445 => D <= "10000010";	-- 0x192D
		when 006446 => D <= "00011000";	-- 0x192E
		when 006447 => D <= "11100010";	-- 0x192F
		when 006448 => D <= "00011101";	-- 0x1930
		when 006449 => D <= "11101101";	-- 0x1931
		when 006450 => D <= "00011010";	-- 0x1932
		when 006451 => D <= "11110011";	-- 0x1933
		when 006452 => D <= "00011010";	-- 0x1934
		when 006453 => D <= "00000011";	-- 0x1935
		when 006454 => D <= "00011011";	-- 0x1936
		when 006455 => D <= "00000011";	-- 0x1937
		when 006456 => D <= "00011011";	-- 0x1938
		when 006457 => D <= "00000011";	-- 0x1939
		when 006458 => D <= "00011011";	-- 0x193A
		when 006459 => D <= "00000011";	-- 0x193B
		when 006460 => D <= "00011011";	-- 0x193C
		when 006461 => D <= "00000011";	-- 0x193D
		when 006462 => D <= "00011011";	-- 0x193E
		when 006463 => D <= "00000011";	-- 0x193F
		when 006464 => D <= "00011011";	-- 0x1940
		when 006465 => D <= "01010101";	-- 0x1941
		when 006466 => D <= "00010111";	-- 0x1942
		when 006467 => D <= "11111000";	-- 0x1943
		when 006468 => D <= "00011010";	-- 0x1944
		when 006469 => D <= "00000011";	-- 0x1945
		when 006470 => D <= "00011011";	-- 0x1946
		when 006471 => D <= "00000011";	-- 0x1947
		when 006472 => D <= "00011011";	-- 0x1948
		when 006473 => D <= "00000011";	-- 0x1949
		when 006474 => D <= "00011011";	-- 0x194A
		when 006475 => D <= "00000011";	-- 0x194B
		when 006476 => D <= "00011011";	-- 0x194C
		when 006477 => D <= "00000011";	-- 0x194D
		when 006478 => D <= "00011011";	-- 0x194E
		when 006479 => D <= "00000011";	-- 0x194F
		when 006480 => D <= "00011011";	-- 0x1950
		when 006481 => D <= "01100010";	-- 0x1951
		when 006482 => D <= "00011011";	-- 0x1952
		when 006483 => D <= "10100000";	-- 0x1953
		when 006484 => D <= "00011010";	-- 0x1954
		when 006485 => D <= "00000110";	-- 0x1955
		when 006486 => D <= "00011100";	-- 0x1956
		when 006487 => D <= "10100100";	-- 0x1957
		when 006488 => D <= "00011011";	-- 0x1958
		when 006489 => D <= "00010001";	-- 0x1959
		when 006490 => D <= "00011100";	-- 0x195A
		when 006491 => D <= "01001001";	-- 0x195B
		when 006492 => D <= "00011101";	-- 0x195C
		when 006493 => D <= "00111110";	-- 0x195D
		when 006494 => D <= "00011101";	-- 0x195E
		when 006495 => D <= "01101110";	-- 0x195F
		when 006496 => D <= "00011101";	-- 0x1960
		when 006497 => D <= "11000100";	-- 0x1961
		when 006498 => D <= "00011101";	-- 0x1962
		when 006499 => D <= "11010100";	-- 0x1963
		when 006500 => D <= "00011101";	-- 0x1964
		when 006501 => D <= "01110110";	-- 0x1965
		when 006502 => D <= "00011101";	-- 0x1966
		when 006503 => D <= "10101001";	-- 0x1967
		when 006504 => D <= "00011100";	-- 0x1968
		when 006505 => D <= "01011011";	-- 0x1969
		when 006506 => D <= "00011100";	-- 0x196A
		when 006507 => D <= "01000110";	-- 0x196B
		when 006508 => D <= "00011100";	-- 0x196C
		when 006509 => D <= "11011011";	-- 0x196D
		when 006510 => D <= "00011101";	-- 0x196E
		when 006511 => D <= "10101111";	-- 0x196F
		when 006512 => D <= "00011010";	-- 0x1970
		when 006513 => D <= "10101010";	-- 0x1971
		when 006514 => D <= "00011010";	-- 0x1972
		when 006515 => D <= "10111110";	-- 0x1973
		when 006516 => D <= "00011010";	-- 0x1974
		when 006517 => D <= "11000101";	-- 0x1975
		when 006518 => D <= "00011010";	-- 0x1976
		when 006519 => D <= "11010101";	-- 0x1977
		when 006520 => D <= "00011011";	-- 0x1978
		when 006521 => D <= "10001111";	-- 0x1979
		when 006522 => D <= "00011011";	-- 0x197A
		when 006523 => D <= "11010101";	-- 0x197B
		when 006524 => D <= "00011010";	-- 0x197C
		when 006525 => D <= "11110110";	-- 0x197D
		when 006526 => D <= "00011001";	-- 0x197E
		when 006527 => D <= "00110111";	-- 0x197F
		when 006528 => D <= "00011100";	-- 0x1980
		when 006529 => D <= "00100011";	-- 0x1981
		when 006530 => D <= "00011100";	-- 0x1982
		when 006531 => D <= "11111100";	-- 0x1983
		when 006532 => D <= "00011001";	-- 0x1984
		when 006533 => D <= "00010111";	-- 0x1985
		when 006534 => D <= "00011100";	-- 0x1986
		when 006535 => D <= "11011011";	-- 0x1987
		when 006536 => D <= "00011010";	-- 0x1988
		when 006537 => D <= "11001110";	-- 0x1989
		when 006538 => D <= "00011010";	-- 0x198A
		when 006539 => D <= "00101011";	-- 0x198B
		when 006540 => D <= "00000000";	-- 0x198C
		when 006541 => D <= "00011000";	-- 0x198D
		when 006542 => D <= "00011101";	-- 0x198E
		when 006543 => D <= "11100100";	-- 0x198F
		when 006544 => D <= "00011000";	-- 0x1990
		when 006545 => D <= "11100100";	-- 0x1991
		when 006546 => D <= "00011001";	-- 0x1992
		when 006547 => D <= "01011010";	-- 0x1993
		when 006548 => D <= "00010101";	-- 0x1994
		when 006549 => D <= "01111111";	-- 0x1995
		when 006550 => D <= "00011010";	-- 0x1996
		when 006551 => D <= "01010001";	-- 0x1997
		when 006552 => D <= "00011010";	-- 0x1998
		when 006553 => D <= "01100011";	-- 0x1999
		when 006554 => D <= "00011010";	-- 0x199A
		when 006555 => D <= "01000101";	-- 0x199B
		when 006556 => D <= "00011010";	-- 0x199C
		when 006557 => D <= "11001101";	-- 0x199D
		when 006558 => D <= "10000101";	-- 0x199E
		when 006559 => D <= "00011011";	-- 0x199F
		when 006560 => D <= "01111000";	-- 0x19A0
		when 006561 => D <= "00110010";	-- 0x19A1
		when 006562 => D <= "00011110";	-- 0x19A2
		when 006563 => D <= "01000000";	-- 0x19A3
		when 006564 => D <= "11011001";	-- 0x19A4
		when 006565 => D <= "11100011";	-- 0x19A5
		when 006566 => D <= "11011001";	-- 0x19A6
		when 006567 => D <= "11101101";	-- 0x19A7
		when 006568 => D <= "01010011";	-- 0x19A8
		when 006569 => D <= "00011100";	-- 0x19A9
		when 006570 => D <= "01000000";	-- 0x19AA
		when 006571 => D <= "11011001";	-- 0x19AB
		when 006572 => D <= "01111110";	-- 0x19AC
		when 006573 => D <= "00100011";	-- 0x19AD
		when 006574 => D <= "11100101";	-- 0x19AE
		when 006575 => D <= "10100111";	-- 0x19AF
		when 006576 => D <= "11110010";	-- 0x19B0
		when 006577 => D <= "11000010";	-- 0x19B1
		when 006578 => D <= "00011001";	-- 0x19B2
		when 006579 => D <= "01010111";	-- 0x19B3
		when 006580 => D <= "11100110";	-- 0x19B4
		when 006581 => D <= "01100000";	-- 0x19B5
		when 006582 => D <= "00001111";	-- 0x19B6
		when 006583 => D <= "00001111";	-- 0x19B7
		when 006584 => D <= "00001111";	-- 0x19B8
		when 006585 => D <= "00001111";	-- 0x19B9
		when 006586 => D <= "11000110";	-- 0x19BA
		when 006587 => D <= "01110010";	-- 0x19BB
		when 006588 => D <= "01101111";	-- 0x19BC
		when 006589 => D <= "01111010";	-- 0x19BD
		when 006590 => D <= "11100110";	-- 0x19BE
		when 006591 => D <= "00011111";	-- 0x19BF
		when 006592 => D <= "00011000";	-- 0x19C0
		when 006593 => D <= "00001110";	-- 0x19C1
		when 006594 => D <= "11111110";	-- 0x19C2
		when 006595 => D <= "00011000";	-- 0x19C3
		when 006596 => D <= "00110000";	-- 0x19C4
		when 006597 => D <= "00001000";	-- 0x19C5
		when 006598 => D <= "11011001";	-- 0x19C6
		when 006599 => D <= "00000001";	-- 0x19C7
		when 006600 => D <= "11111011";	-- 0x19C8
		when 006601 => D <= "11111111";	-- 0x19C9
		when 006602 => D <= "01010100";	-- 0x19CA
		when 006603 => D <= "01011101";	-- 0x19CB
		when 006604 => D <= "00001001";	-- 0x19CC
		when 006605 => D <= "11011001";	-- 0x19CD
		when 006606 => D <= "00000111";	-- 0x19CE
		when 006607 => D <= "01101111";	-- 0x19CF
		when 006608 => D <= "00010001";	-- 0x19D0
		when 006609 => D <= "00100011";	-- 0x19D1
		when 006610 => D <= "00011001";	-- 0x19D2
		when 006611 => D <= "00100110";	-- 0x19D3
		when 006612 => D <= "00000000";	-- 0x19D4
		when 006613 => D <= "00011001";	-- 0x19D5
		when 006614 => D <= "01011110";	-- 0x19D6
		when 006615 => D <= "00100011";	-- 0x19D7
		when 006616 => D <= "01010110";	-- 0x19D8
		when 006617 => D <= "00100001";	-- 0x19D9
		when 006618 => D <= "10100111";	-- 0x19DA
		when 006619 => D <= "00011001";	-- 0x19DB
		when 006620 => D <= "11100011";	-- 0x19DC
		when 006621 => D <= "11010101";	-- 0x19DD
		when 006622 => D <= "11011001";	-- 0x19DE
		when 006623 => D <= "11101101";	-- 0x19DF
		when 006624 => D <= "01001011";	-- 0x19E0
		when 006625 => D <= "00011101";	-- 0x19E1
		when 006626 => D <= "01000000";	-- 0x19E2
		when 006627 => D <= "11001001";	-- 0x19E3
		when 006628 => D <= "11110001";	-- 0x19E4
		when 006629 => D <= "00111010";	-- 0x19E5
		when 006630 => D <= "00011110";	-- 0x19E6
		when 006631 => D <= "01000000";	-- 0x19E7
		when 006632 => D <= "11011001";	-- 0x19E8
		when 006633 => D <= "00011000";	-- 0x19E9
		when 006634 => D <= "11000011";	-- 0x19EA
		when 006635 => D <= "11010101";	-- 0x19EB
		when 006636 => D <= "11100101";	-- 0x19EC
		when 006637 => D <= "00000001";	-- 0x19ED
		when 006638 => D <= "00000101";	-- 0x19EE
		when 006639 => D <= "00000000";	-- 0x19EF
		when 006640 => D <= "11001101";	-- 0x19F0
		when 006641 => D <= "11000101";	-- 0x19F1
		when 006642 => D <= "00001110";	-- 0x19F2
		when 006643 => D <= "11100001";	-- 0x19F3
		when 006644 => D <= "11010001";	-- 0x19F4
		when 006645 => D <= "11001001";	-- 0x19F5
		when 006646 => D <= "11001101";	-- 0x19F6
		when 006647 => D <= "11101011";	-- 0x19F7
		when 006648 => D <= "00011001";	-- 0x19F8
		when 006649 => D <= "11101101";	-- 0x19F9
		when 006650 => D <= "10110000";	-- 0x19FA
		when 006651 => D <= "11001001";	-- 0x19FB
		when 006652 => D <= "01100010";	-- 0x19FC
		when 006653 => D <= "01101011";	-- 0x19FD
		when 006654 => D <= "11001101";	-- 0x19FE
		when 006655 => D <= "11101011";	-- 0x19FF
		when 006656 => D <= "00011001";	-- 0x1A00
		when 006657 => D <= "11011001";	-- 0x1A01
		when 006658 => D <= "11100101";	-- 0x1A02
		when 006659 => D <= "11011001";	-- 0x1A03
		when 006660 => D <= "11100011";	-- 0x1A04
		when 006661 => D <= "11000101";	-- 0x1A05
		when 006662 => D <= "01111110";	-- 0x1A06
		when 006663 => D <= "11100110";	-- 0x1A07
		when 006664 => D <= "11000000";	-- 0x1A08
		when 006665 => D <= "00000111";	-- 0x1A09
		when 006666 => D <= "00000111";	-- 0x1A0A
		when 006667 => D <= "01001111";	-- 0x1A0B
		when 006668 => D <= "00001100";	-- 0x1A0C
		when 006669 => D <= "01111110";	-- 0x1A0D
		when 006670 => D <= "11100110";	-- 0x1A0E
		when 006671 => D <= "00111111";	-- 0x1A0F
		when 006672 => D <= "00100000";	-- 0x1A10
		when 006673 => D <= "00000010";	-- 0x1A11
		when 006674 => D <= "00100011";	-- 0x1A12
		when 006675 => D <= "01111110";	-- 0x1A13
		when 006676 => D <= "11000110";	-- 0x1A14
		when 006677 => D <= "01010000";	-- 0x1A15
		when 006678 => D <= "00010010";	-- 0x1A16
		when 006679 => D <= "00111110";	-- 0x1A17
		when 006680 => D <= "00000101";	-- 0x1A18
		when 006681 => D <= "10010001";	-- 0x1A19
		when 006682 => D <= "00100011";	-- 0x1A1A
		when 006683 => D <= "00010011";	-- 0x1A1B
		when 006684 => D <= "00000110";	-- 0x1A1C
		when 006685 => D <= "00000000";	-- 0x1A1D
		when 006686 => D <= "11101101";	-- 0x1A1E
		when 006687 => D <= "10110000";	-- 0x1A1F
		when 006688 => D <= "11000001";	-- 0x1A20
		when 006689 => D <= "11100011";	-- 0x1A21
		when 006690 => D <= "11011001";	-- 0x1A22
		when 006691 => D <= "11100001";	-- 0x1A23
		when 006692 => D <= "11011001";	-- 0x1A24
		when 006693 => D <= "01000111";	-- 0x1A25
		when 006694 => D <= "10101111";	-- 0x1A26
		when 006695 => D <= "00000101";	-- 0x1A27
		when 006696 => D <= "11001000";	-- 0x1A28
		when 006697 => D <= "00010010";	-- 0x1A29
		when 006698 => D <= "00010011";	-- 0x1A2A
		when 006699 => D <= "00011000";	-- 0x1A2B
		when 006700 => D <= "11111010";	-- 0x1A2C
		when 006701 => D <= "10100111";	-- 0x1A2D
		when 006702 => D <= "11001000";	-- 0x1A2E
		when 006703 => D <= "11110101";	-- 0x1A2F
		when 006704 => D <= "11010101";	-- 0x1A30
		when 006705 => D <= "00010001";	-- 0x1A31
		when 006706 => D <= "00000000";	-- 0x1A32
		when 006707 => D <= "00000000";	-- 0x1A33
		when 006708 => D <= "11001101";	-- 0x1A34
		when 006709 => D <= "11111110";	-- 0x1A35
		when 006710 => D <= "00011001";	-- 0x1A36
		when 006711 => D <= "11010001";	-- 0x1A37
		when 006712 => D <= "11110001";	-- 0x1A38
		when 006713 => D <= "00111101";	-- 0x1A39
		when 006714 => D <= "00011000";	-- 0x1A3A
		when 006715 => D <= "11110010";	-- 0x1A3B
		when 006716 => D <= "01001111";	-- 0x1A3C
		when 006717 => D <= "00000111";	-- 0x1A3D
		when 006718 => D <= "00000111";	-- 0x1A3E
		when 006719 => D <= "10000001";	-- 0x1A3F
		when 006720 => D <= "01001111";	-- 0x1A40
		when 006721 => D <= "00000110";	-- 0x1A41
		when 006722 => D <= "00000000";	-- 0x1A42
		when 006723 => D <= "00001001";	-- 0x1A43
		when 006724 => D <= "11001001";	-- 0x1A44
		when 006725 => D <= "11010101";	-- 0x1A45
		when 006726 => D <= "00101010";	-- 0x1A46
		when 006727 => D <= "00011111";	-- 0x1A47
		when 006728 => D <= "01000000";	-- 0x1A48
		when 006729 => D <= "11001101";	-- 0x1A49
		when 006730 => D <= "00111100";	-- 0x1A4A
		when 006731 => D <= "00011010";	-- 0x1A4B
		when 006732 => D <= "11001101";	-- 0x1A4C
		when 006733 => D <= "11110110";	-- 0x1A4D
		when 006734 => D <= "00011001";	-- 0x1A4E
		when 006735 => D <= "11100001";	-- 0x1A4F
		when 006736 => D <= "11001001";	-- 0x1A50
		when 006737 => D <= "01100010";	-- 0x1A51
		when 006738 => D <= "01101011";	-- 0x1A52
		when 006739 => D <= "11011001";	-- 0x1A53
		when 006740 => D <= "11100101";	-- 0x1A54
		when 006741 => D <= "00100001";	-- 0x1A55
		when 006742 => D <= "00010101";	-- 0x1A56
		when 006743 => D <= "00011001";	-- 0x1A57
		when 006744 => D <= "11011001";	-- 0x1A58
		when 006745 => D <= "11001101";	-- 0x1A59
		when 006746 => D <= "00101101";	-- 0x1A5A
		when 006747 => D <= "00011010";	-- 0x1A5B
		when 006748 => D <= "11001101";	-- 0x1A5C
		when 006749 => D <= "11111110";	-- 0x1A5D
		when 006750 => D <= "00011001";	-- 0x1A5E
		when 006751 => D <= "11011001";	-- 0x1A5F
		when 006752 => D <= "11100001";	-- 0x1A60
		when 006753 => D <= "11011001";	-- 0x1A61
		when 006754 => D <= "11001001";	-- 0x1A62
		when 006755 => D <= "11100101";	-- 0x1A63
		when 006756 => D <= "11101011";	-- 0x1A64
		when 006757 => D <= "00101010";	-- 0x1A65
		when 006758 => D <= "00011111";	-- 0x1A66
		when 006759 => D <= "01000000";	-- 0x1A67
		when 006760 => D <= "11001101";	-- 0x1A68
		when 006761 => D <= "00111100";	-- 0x1A69
		when 006762 => D <= "00011010";	-- 0x1A6A
		when 006763 => D <= "11101011";	-- 0x1A6B
		when 006764 => D <= "11001101";	-- 0x1A6C
		when 006765 => D <= "11110110";	-- 0x1A6D
		when 006766 => D <= "00011001";	-- 0x1A6E
		when 006767 => D <= "11101011";	-- 0x1A6F
		when 006768 => D <= "11100001";	-- 0x1A70
		when 006769 => D <= "11001001";	-- 0x1A71
		when 006770 => D <= "00000110";	-- 0x1A72
		when 006771 => D <= "00000101";	-- 0x1A73
		when 006772 => D <= "00011010";	-- 0x1A74
		when 006773 => D <= "01001110";	-- 0x1A75
		when 006774 => D <= "11101011";	-- 0x1A76
		when 006775 => D <= "00010010";	-- 0x1A77
		when 006776 => D <= "01110001";	-- 0x1A78
		when 006777 => D <= "00100011";	-- 0x1A79
		when 006778 => D <= "00010011";	-- 0x1A7A
		when 006779 => D <= "00010000";	-- 0x1A7B
		when 006780 => D <= "11110111";	-- 0x1A7C
		when 006781 => D <= "11101011";	-- 0x1A7D
		when 006782 => D <= "11001001";	-- 0x1A7E
		when 006783 => D <= "01000111";	-- 0x1A7F
		when 006784 => D <= "11001101";	-- 0x1A80
		when 006785 => D <= "10100000";	-- 0x1A81
		when 006786 => D <= "00011001";	-- 0x1A82
		when 006787 => D <= "00101101";	-- 0x1A83
		when 006788 => D <= "00001111";	-- 0x1A84
		when 006789 => D <= "11000000";	-- 0x1A85
		when 006790 => D <= "00000010";	-- 0x1A86
		when 006791 => D <= "10100000";	-- 0x1A87
		when 006792 => D <= "11000010";	-- 0x1A88
		when 006793 => D <= "00101101";	-- 0x1A89
		when 006794 => D <= "11100000";	-- 0x1A8A
		when 006795 => D <= "00000100";	-- 0x1A8B
		when 006796 => D <= "11100010";	-- 0x1A8C
		when 006797 => D <= "11000001";	-- 0x1A8D
		when 006798 => D <= "00000011";	-- 0x1A8E
		when 006799 => D <= "00110100";	-- 0x1A8F
		when 006800 => D <= "11001101";	-- 0x1A90
		when 006801 => D <= "11111100";	-- 0x1A91
		when 006802 => D <= "00011001";	-- 0x1A92
		when 006803 => D <= "11001101";	-- 0x1A93
		when 006804 => D <= "10100100";	-- 0x1A94
		when 006805 => D <= "00011001";	-- 0x1A95
		when 006806 => D <= "00001111";	-- 0x1A96
		when 006807 => D <= "00000001";	-- 0x1A97
		when 006808 => D <= "11000010";	-- 0x1A98
		when 006809 => D <= "00000010";	-- 0x1A99
		when 006810 => D <= "00110001";	-- 0x1A9A
		when 006811 => D <= "11101110";	-- 0x1A9B
		when 006812 => D <= "11100001";	-- 0x1A9C
		when 006813 => D <= "00000011";	-- 0x1A9D
		when 006814 => D <= "00110100";	-- 0x1A9E
		when 006815 => D <= "11001001";	-- 0x1A9F
		when 006816 => D <= "01111110";	-- 0x1AA0
		when 006817 => D <= "10100111";	-- 0x1AA1
		when 006818 => D <= "11001000";	-- 0x1AA2
		when 006819 => D <= "00100011";	-- 0x1AA3
		when 006820 => D <= "01111110";	-- 0x1AA4
		when 006821 => D <= "11101110";	-- 0x1AA5
		when 006822 => D <= "10000000";	-- 0x1AA6
		when 006823 => D <= "01110111";	-- 0x1AA7
		when 006824 => D <= "00101011";	-- 0x1AA8
		when 006825 => D <= "11001001";	-- 0x1AA9
		when 006826 => D <= "00100011";	-- 0x1AAA
		when 006827 => D <= "11001011";	-- 0x1AAB
		when 006828 => D <= "10111110";	-- 0x1AAC
		when 006829 => D <= "00101011";	-- 0x1AAD
		when 006830 => D <= "11001001";	-- 0x1AAE
		when 006831 => D <= "00100011";	-- 0x1AAF
		when 006832 => D <= "01111110";	-- 0x1AB0
		when 006833 => D <= "00101011";	-- 0x1AB1
		when 006834 => D <= "00110101";	-- 0x1AB2
		when 006835 => D <= "00110100";	-- 0x1AB3
		when 006836 => D <= "00110111";	-- 0x1AB4
		when 006837 => D <= "11000100";	-- 0x1AB5
		when 006838 => D <= "11100000";	-- 0x1AB6
		when 006839 => D <= "00011010";	-- 0x1AB7
		when 006840 => D <= "00100011";	-- 0x1AB8
		when 006841 => D <= "00000111";	-- 0x1AB9
		when 006842 => D <= "11001011";	-- 0x1ABA
		when 006843 => D <= "00011110";	-- 0x1ABB
		when 006844 => D <= "00101011";	-- 0x1ABC
		when 006845 => D <= "11001001";	-- 0x1ABD
		when 006846 => D <= "11001101";	-- 0x1ABE
		when 006847 => D <= "10100111";	-- 0x1ABF
		when 006848 => D <= "00001110";	-- 0x1AC0
		when 006849 => D <= "00001010";	-- 0x1AC1
		when 006850 => D <= "11000011";	-- 0x1AC2
		when 006851 => D <= "00011101";	-- 0x1AC3
		when 006852 => D <= "00010101";	-- 0x1AC4
		when 006853 => D <= "11001101";	-- 0x1AC5
		when 006854 => D <= "10100111";	-- 0x1AC6
		when 006855 => D <= "00001110";	-- 0x1AC7
		when 006856 => D <= "00100001";	-- 0x1AC8
		when 006857 => D <= "00100000";	-- 0x1AC9
		when 006858 => D <= "00010101";	-- 0x1ACA
		when 006859 => D <= "11100101";	-- 0x1ACB
		when 006860 => D <= "11000101";	-- 0x1ACC
		when 006861 => D <= "11001001";	-- 0x1ACD
		when 006862 => D <= "01111110";	-- 0x1ACE
		when 006863 => D <= "10100111";	-- 0x1ACF
		when 006864 => D <= "11001000";	-- 0x1AD0
		when 006865 => D <= "00111110";	-- 0x1AD1
		when 006866 => D <= "11111111";	-- 0x1AD2
		when 006867 => D <= "00011000";	-- 0x1AD3
		when 006868 => D <= "00000111";	-- 0x1AD4
		when 006869 => D <= "01111110";	-- 0x1AD5
		when 006870 => D <= "11101101";	-- 0x1AD6
		when 006871 => D <= "01000100";	-- 0x1AD7
		when 006872 => D <= "00111111";	-- 0x1AD8
		when 006873 => D <= "00011000";	-- 0x1AD9
		when 006874 => D <= "00000101";	-- 0x1ADA
		when 006875 => D <= "10101111";	-- 0x1ADB
		when 006876 => D <= "00100011";	-- 0x1ADC
		when 006877 => D <= "10101110";	-- 0x1ADD
		when 006878 => D <= "00101011";	-- 0x1ADE
		when 006879 => D <= "00000111";	-- 0x1ADF
		when 006880 => D <= "11100101";	-- 0x1AE0
		when 006881 => D <= "00000110";	-- 0x1AE1
		when 006882 => D <= "00000101";	-- 0x1AE2
		when 006883 => D <= "00110110";	-- 0x1AE3
		when 006884 => D <= "00000000";	-- 0x1AE4
		when 006885 => D <= "00100011";	-- 0x1AE5
		when 006886 => D <= "00010000";	-- 0x1AE6
		when 006887 => D <= "11111011";	-- 0x1AE7
		when 006888 => D <= "11100001";	-- 0x1AE8
		when 006889 => D <= "11010000";	-- 0x1AE9
		when 006890 => D <= "00110110";	-- 0x1AEA
		when 006891 => D <= "10000001";	-- 0x1AEB
		when 006892 => D <= "11001001";	-- 0x1AEC
		when 006893 => D <= "00011010";	-- 0x1AED
		when 006894 => D <= "10100111";	-- 0x1AEE
		when 006895 => D <= "11001000";	-- 0x1AEF
		when 006896 => D <= "00110111";	-- 0x1AF0
		when 006897 => D <= "00011000";	-- 0x1AF1
		when 006898 => D <= "11101101";	-- 0x1AF2
		when 006899 => D <= "00011010";	-- 0x1AF3
		when 006900 => D <= "10100111";	-- 0x1AF4
		when 006901 => D <= "11000000";	-- 0x1AF5
		when 006902 => D <= "00011000";	-- 0x1AF6
		when 006903 => D <= "11101000";	-- 0x1AF7
		when 006904 => D <= "00011010";	-- 0x1AF8
		when 006905 => D <= "10100111";	-- 0x1AF9
		when 006906 => D <= "11000000";	-- 0x1AFA
		when 006907 => D <= "11010101";	-- 0x1AFB
		when 006908 => D <= "00011011";	-- 0x1AFC
		when 006909 => D <= "10101111";	-- 0x1AFD
		when 006910 => D <= "00010010";	-- 0x1AFE
		when 006911 => D <= "00011011";	-- 0x1AFF
		when 006912 => D <= "00010010";	-- 0x1B00
		when 006913 => D <= "11010001";	-- 0x1B01
		when 006914 => D <= "11001001";	-- 0x1B02
		when 006915 => D <= "01111000";	-- 0x1B03
		when 006916 => D <= "11010110";	-- 0x1B04
		when 006917 => D <= "00001000";	-- 0x1B05
		when 006918 => D <= "11001011";	-- 0x1B06
		when 006919 => D <= "01010111";	-- 0x1B07
		when 006920 => D <= "00100000";	-- 0x1B08
		when 006921 => D <= "00000001";	-- 0x1B09
		when 006922 => D <= "00111101";	-- 0x1B0A
		when 006923 => D <= "00001111";	-- 0x1B0B
		when 006924 => D <= "00110000";	-- 0x1B0C
		when 006925 => D <= "00001000";	-- 0x1B0D
		when 006926 => D <= "11110101";	-- 0x1B0E
		when 006927 => D <= "11100101";	-- 0x1B0F
		when 006928 => D <= "11001101";	-- 0x1B10
		when 006929 => D <= "01110010";	-- 0x1B11
		when 006930 => D <= "00011010";	-- 0x1B12
		when 006931 => D <= "11010001";	-- 0x1B13
		when 006932 => D <= "11101011";	-- 0x1B14
		when 006933 => D <= "11110001";	-- 0x1B15
		when 006934 => D <= "11001011";	-- 0x1B16
		when 006935 => D <= "01010111";	-- 0x1B17
		when 006936 => D <= "00100000";	-- 0x1B18
		when 006937 => D <= "00000111";	-- 0x1B19
		when 006938 => D <= "00001111";	-- 0x1B1A
		when 006939 => D <= "11110101";	-- 0x1B1B
		when 006940 => D <= "11001101";	-- 0x1B1C
		when 006941 => D <= "01001100";	-- 0x1B1D
		when 006942 => D <= "00010111";	-- 0x1B1E
		when 006943 => D <= "00011000";	-- 0x1B1F
		when 006944 => D <= "00110011";	-- 0x1B20
		when 006945 => D <= "00001111";	-- 0x1B21
		when 006946 => D <= "11110101";	-- 0x1B22
		when 006947 => D <= "11001101";	-- 0x1B23
		when 006948 => D <= "11111000";	-- 0x1B24
		when 006949 => D <= "00010011";	-- 0x1B25
		when 006950 => D <= "11010101";	-- 0x1B26
		when 006951 => D <= "11000101";	-- 0x1B27
		when 006952 => D <= "11001101";	-- 0x1B28
		when 006953 => D <= "11111000";	-- 0x1B29
		when 006954 => D <= "00010011";	-- 0x1B2A
		when 006955 => D <= "11100001";	-- 0x1B2B
		when 006956 => D <= "01111100";	-- 0x1B2C
		when 006957 => D <= "10110101";	-- 0x1B2D
		when 006958 => D <= "11100011";	-- 0x1B2E
		when 006959 => D <= "01111000";	-- 0x1B2F
		when 006960 => D <= "00100000";	-- 0x1B30
		when 006961 => D <= "00001011";	-- 0x1B31
		when 006962 => D <= "10110001";	-- 0x1B32
		when 006963 => D <= "11000001";	-- 0x1B33
		when 006964 => D <= "00101000";	-- 0x1B34
		when 006965 => D <= "00000100";	-- 0x1B35
		when 006966 => D <= "11110001";	-- 0x1B36
		when 006967 => D <= "00111111";	-- 0x1B37
		when 006968 => D <= "00011000";	-- 0x1B38
		when 006969 => D <= "00010110";	-- 0x1B39
		when 006970 => D <= "11110001";	-- 0x1B3A
		when 006971 => D <= "00011000";	-- 0x1B3B
		when 006972 => D <= "00010011";	-- 0x1B3C
		when 006973 => D <= "10110001";	-- 0x1B3D
		when 006974 => D <= "00101000";	-- 0x1B3E
		when 006975 => D <= "00001101";	-- 0x1B3F
		when 006976 => D <= "00011010";	-- 0x1B40
		when 006977 => D <= "10010110";	-- 0x1B41
		when 006978 => D <= "00111000";	-- 0x1B42
		when 006979 => D <= "00001001";	-- 0x1B43
		when 006980 => D <= "00100000";	-- 0x1B44
		when 006981 => D <= "11101101";	-- 0x1B45
		when 006982 => D <= "00001011";	-- 0x1B46
		when 006983 => D <= "00010011";	-- 0x1B47
		when 006984 => D <= "00100011";	-- 0x1B48
		when 006985 => D <= "11100011";	-- 0x1B49
		when 006986 => D <= "00101011";	-- 0x1B4A
		when 006987 => D <= "00011000";	-- 0x1B4B
		when 006988 => D <= "11011111";	-- 0x1B4C
		when 006989 => D <= "11000001";	-- 0x1B4D
		when 006990 => D <= "11110001";	-- 0x1B4E
		when 006991 => D <= "10100111";	-- 0x1B4F
		when 006992 => D <= "11110101";	-- 0x1B50
		when 006993 => D <= "11101111";	-- 0x1B51
		when 006994 => D <= "10100000";	-- 0x1B52
		when 006995 => D <= "00110100";	-- 0x1B53
		when 006996 => D <= "11110001";	-- 0x1B54
		when 006997 => D <= "11110101";	-- 0x1B55
		when 006998 => D <= "11011100";	-- 0x1B56
		when 006999 => D <= "11010101";	-- 0x1B57
		when 007000 => D <= "00011010";	-- 0x1B58
		when 007001 => D <= "11001101";	-- 0x1B59
		when 007002 => D <= "11001110";	-- 0x1B5A
		when 007003 => D <= "00011010";	-- 0x1B5B
		when 007004 => D <= "11110001";	-- 0x1B5C
		when 007005 => D <= "00001111";	-- 0x1B5D
		when 007006 => D <= "11010100";	-- 0x1B5E
		when 007007 => D <= "11010101";	-- 0x1B5F
		when 007008 => D <= "00011010";	-- 0x1B60
		when 007009 => D <= "11001001";	-- 0x1B61
		when 007010 => D <= "11001101";	-- 0x1B62
		when 007011 => D <= "11111000";	-- 0x1B63
		when 007012 => D <= "00010011";	-- 0x1B64
		when 007013 => D <= "11010101";	-- 0x1B65
		when 007014 => D <= "11000101";	-- 0x1B66
		when 007015 => D <= "11001101";	-- 0x1B67
		when 007016 => D <= "11111000";	-- 0x1B68
		when 007017 => D <= "00010011";	-- 0x1B69
		when 007018 => D <= "11100001";	-- 0x1B6A
		when 007019 => D <= "11100101";	-- 0x1B6B
		when 007020 => D <= "11010101";	-- 0x1B6C
		when 007021 => D <= "11000101";	-- 0x1B6D
		when 007022 => D <= "00001001";	-- 0x1B6E
		when 007023 => D <= "01000100";	-- 0x1B6F
		when 007024 => D <= "01001101";	-- 0x1B70
		when 007025 => D <= "11110111";	-- 0x1B71
		when 007026 => D <= "11001101";	-- 0x1B72
		when 007027 => D <= "11000011";	-- 0x1B73
		when 007028 => D <= "00010010";	-- 0x1B74
		when 007029 => D <= "11000001";	-- 0x1B75
		when 007030 => D <= "11100001";	-- 0x1B76
		when 007031 => D <= "01111000";	-- 0x1B77
		when 007032 => D <= "10110001";	-- 0x1B78
		when 007033 => D <= "00101000";	-- 0x1B79
		when 007034 => D <= "00000010";	-- 0x1B7A
		when 007035 => D <= "11101101";	-- 0x1B7B
		when 007036 => D <= "10110000";	-- 0x1B7C
		when 007037 => D <= "11000001";	-- 0x1B7D
		when 007038 => D <= "11100001";	-- 0x1B7E
		when 007039 => D <= "01111000";	-- 0x1B7F
		when 007040 => D <= "10110001";	-- 0x1B80
		when 007041 => D <= "00101000";	-- 0x1B81
		when 007042 => D <= "00000010";	-- 0x1B82
		when 007043 => D <= "11101101";	-- 0x1B83
		when 007044 => D <= "10110000";	-- 0x1B84
		when 007045 => D <= "00101010";	-- 0x1B85
		when 007046 => D <= "00011100";	-- 0x1B86
		when 007047 => D <= "01000000";	-- 0x1B87
		when 007048 => D <= "00010001";	-- 0x1B88
		when 007049 => D <= "11111011";	-- 0x1B89
		when 007050 => D <= "11111111";	-- 0x1B8A
		when 007051 => D <= "11100101";	-- 0x1B8B
		when 007052 => D <= "00011001";	-- 0x1B8C
		when 007053 => D <= "11010001";	-- 0x1B8D
		when 007054 => D <= "11001001";	-- 0x1B8E
		when 007055 => D <= "11001101";	-- 0x1B8F
		when 007056 => D <= "11001101";	-- 0x1B90
		when 007057 => D <= "00010101";	-- 0x1B91
		when 007058 => D <= "00111000";	-- 0x1B92
		when 007059 => D <= "00001110";	-- 0x1B93
		when 007060 => D <= "00100000";	-- 0x1B94
		when 007061 => D <= "00001100";	-- 0x1B95
		when 007062 => D <= "11110101";	-- 0x1B96
		when 007063 => D <= "00000001";	-- 0x1B97
		when 007064 => D <= "00000001";	-- 0x1B98
		when 007065 => D <= "00000000";	-- 0x1B99
		when 007066 => D <= "11110111";	-- 0x1B9A
		when 007067 => D <= "11110001";	-- 0x1B9B
		when 007068 => D <= "00010010";	-- 0x1B9C
		when 007069 => D <= "11001101";	-- 0x1B9D
		when 007070 => D <= "11000011";	-- 0x1B9E
		when 007071 => D <= "00010010";	-- 0x1B9F
		when 007072 => D <= "11101011";	-- 0x1BA0
		when 007073 => D <= "11001001";	-- 0x1BA1
		when 007074 => D <= "11001111";	-- 0x1BA2
		when 007075 => D <= "00001010";	-- 0x1BA3
		when 007076 => D <= "00101010";	-- 0x1BA4
		when 007077 => D <= "00010110";	-- 0x1BA5
		when 007078 => D <= "01000000";	-- 0x1BA6
		when 007079 => D <= "11100101";	-- 0x1BA7
		when 007080 => D <= "11001101";	-- 0x1BA8
		when 007081 => D <= "11111000";	-- 0x1BA9
		when 007082 => D <= "00010011";	-- 0x1BAA
		when 007083 => D <= "11010101";	-- 0x1BAB
		when 007084 => D <= "00000011";	-- 0x1BAC
		when 007085 => D <= "11110111";	-- 0x1BAD
		when 007086 => D <= "11100001";	-- 0x1BAE
		when 007087 => D <= "11101101";	-- 0x1BAF
		when 007088 => D <= "01010011";	-- 0x1BB0
		when 007089 => D <= "00010110";	-- 0x1BB1
		when 007090 => D <= "01000000";	-- 0x1BB2
		when 007091 => D <= "11010101";	-- 0x1BB3
		when 007092 => D <= "11101101";	-- 0x1BB4
		when 007093 => D <= "10110000";	-- 0x1BB5
		when 007094 => D <= "11101011";	-- 0x1BB6
		when 007095 => D <= "00101011";	-- 0x1BB7
		when 007096 => D <= "00110110";	-- 0x1BB8
		when 007097 => D <= "01110110";	-- 0x1BB9
		when 007098 => D <= "11111101";	-- 0x1BBA
		when 007099 => D <= "11001011";	-- 0x1BBB
		when 007100 => D <= "00000001";	-- 0x1BBC
		when 007101 => D <= "10111110";	-- 0x1BBD
		when 007102 => D <= "11001101";	-- 0x1BBE
		when 007103 => D <= "10010010";	-- 0x1BBF
		when 007104 => D <= "00001101";	-- 0x1BC0
		when 007105 => D <= "11001101";	-- 0x1BC1
		when 007106 => D <= "00100010";	-- 0x1BC2
		when 007107 => D <= "00001101";	-- 0x1BC3
		when 007108 => D <= "11100001";	-- 0x1BC4
		when 007109 => D <= "00100010";	-- 0x1BC5
		when 007110 => D <= "00010110";	-- 0x1BC6
		when 007111 => D <= "01000000";	-- 0x1BC7
		when 007112 => D <= "11111101";	-- 0x1BC8
		when 007113 => D <= "11001011";	-- 0x1BC9
		when 007114 => D <= "00000001";	-- 0x1BCA
		when 007115 => D <= "11111110";	-- 0x1BCB
		when 007116 => D <= "11001101";	-- 0x1BCC
		when 007117 => D <= "01010101";	-- 0x1BCD
		when 007118 => D <= "00001111";	-- 0x1BCE
		when 007119 => D <= "11100001";	-- 0x1BCF
		when 007120 => D <= "00100010";	-- 0x1BD0
		when 007121 => D <= "00010110";	-- 0x1BD1
		when 007122 => D <= "01000000";	-- 0x1BD2
		when 007123 => D <= "00011000";	-- 0x1BD3
		when 007124 => D <= "10110000";	-- 0x1BD4
		when 007125 => D <= "00000001";	-- 0x1BD5
		when 007126 => D <= "00000001";	-- 0x1BD6
		when 007127 => D <= "00000000";	-- 0x1BD7
		when 007128 => D <= "11110111";	-- 0x1BD8
		when 007129 => D <= "00110110";	-- 0x1BD9
		when 007130 => D <= "01110110";	-- 0x1BDA
		when 007131 => D <= "00101010";	-- 0x1BDB
		when 007132 => D <= "00111001";	-- 0x1BDC
		when 007133 => D <= "01000000";	-- 0x1BDD
		when 007134 => D <= "11100101";	-- 0x1BDE
		when 007135 => D <= "00101110";	-- 0x1BDF
		when 007136 => D <= "11111111";	-- 0x1BE0
		when 007137 => D <= "00100010";	-- 0x1BE1
		when 007138 => D <= "00111001";	-- 0x1BE2
		when 007139 => D <= "01000000";	-- 0x1BE3
		when 007140 => D <= "00101010";	-- 0x1BE4
		when 007141 => D <= "00001110";	-- 0x1BE5
		when 007142 => D <= "01000000";	-- 0x1BE6
		when 007143 => D <= "11100101";	-- 0x1BE7
		when 007144 => D <= "11101101";	-- 0x1BE8
		when 007145 => D <= "01010011";	-- 0x1BE9
		when 007146 => D <= "00001110";	-- 0x1BEA
		when 007147 => D <= "01000000";	-- 0x1BEB
		when 007148 => D <= "11010101";	-- 0x1BEC
		when 007149 => D <= "11001101";	-- 0x1BED
		when 007150 => D <= "11011011";	-- 0x1BEE
		when 007151 => D <= "00010101";	-- 0x1BEF
		when 007152 => D <= "11010001";	-- 0x1BF0
		when 007153 => D <= "00101010";	-- 0x1BF1
		when 007154 => D <= "00001110";	-- 0x1BF2
		when 007155 => D <= "01000000";	-- 0x1BF3
		when 007156 => D <= "10100111";	-- 0x1BF4
		when 007157 => D <= "11101101";	-- 0x1BF5
		when 007158 => D <= "01010010";	-- 0x1BF6
		when 007159 => D <= "01000100";	-- 0x1BF7
		when 007160 => D <= "01001101";	-- 0x1BF8
		when 007161 => D <= "11100001";	-- 0x1BF9
		when 007162 => D <= "00100010";	-- 0x1BFA
		when 007163 => D <= "00001110";	-- 0x1BFB
		when 007164 => D <= "01000000";	-- 0x1BFC
		when 007165 => D <= "11100001";	-- 0x1BFD
		when 007166 => D <= "00100010";	-- 0x1BFE
		when 007167 => D <= "00111001";	-- 0x1BFF
		when 007168 => D <= "01000000";	-- 0x1C00
		when 007169 => D <= "11001101";	-- 0x1C01
		when 007170 => D <= "11000011";	-- 0x1C02
		when 007171 => D <= "00010010";	-- 0x1C03
		when 007172 => D <= "11101011";	-- 0x1C04
		when 007173 => D <= "11001001";	-- 0x1C05
		when 007174 => D <= "11001101";	-- 0x1C06
		when 007175 => D <= "11111000";	-- 0x1C07
		when 007176 => D <= "00010011";	-- 0x1C08
		when 007177 => D <= "01111000";	-- 0x1C09
		when 007178 => D <= "10110001";	-- 0x1C0A
		when 007179 => D <= "00101000";	-- 0x1C0B
		when 007180 => D <= "00000001";	-- 0x1C0C
		when 007181 => D <= "00011010";	-- 0x1C0D
		when 007182 => D <= "11000011";	-- 0x1C0E
		when 007183 => D <= "00011101";	-- 0x1C0F
		when 007184 => D <= "00010101";	-- 0x1C10
		when 007185 => D <= "11001101";	-- 0x1C11
		when 007186 => D <= "11111000";	-- 0x1C12
		when 007187 => D <= "00010011";	-- 0x1C13
		when 007188 => D <= "11000011";	-- 0x1C14
		when 007189 => D <= "00100000";	-- 0x1C15
		when 007190 => D <= "00010101";	-- 0x1C16
		when 007191 => D <= "11011001";	-- 0x1C17
		when 007192 => D <= "11100101";	-- 0x1C18
		when 007193 => D <= "00100001";	-- 0x1C19
		when 007194 => D <= "00011110";	-- 0x1C1A
		when 007195 => D <= "01000000";	-- 0x1C1B
		when 007196 => D <= "00110101";	-- 0x1C1C
		when 007197 => D <= "11100001";	-- 0x1C1D
		when 007198 => D <= "00100000";	-- 0x1C1E
		when 007199 => D <= "00000100";	-- 0x1C1F
		when 007200 => D <= "00100011";	-- 0x1C20
		when 007201 => D <= "11011001";	-- 0x1C21
		when 007202 => D <= "11001001";	-- 0x1C22
		when 007203 => D <= "11011001";	-- 0x1C23
		when 007204 => D <= "01011110";	-- 0x1C24
		when 007205 => D <= "10101111";	-- 0x1C25
		when 007206 => D <= "11001011";	-- 0x1C26
		when 007207 => D <= "01111011";	-- 0x1C27
		when 007208 => D <= "00101000";	-- 0x1C28
		when 007209 => D <= "00000001";	-- 0x1C29
		when 007210 => D <= "00101111";	-- 0x1C2A
		when 007211 => D <= "01010111";	-- 0x1C2B
		when 007212 => D <= "00011001";	-- 0x1C2C
		when 007213 => D <= "11011001";	-- 0x1C2D
		when 007214 => D <= "11001001";	-- 0x1C2E
		when 007215 => D <= "00011010";	-- 0x1C2F
		when 007216 => D <= "10100111";	-- 0x1C30
		when 007217 => D <= "00100000";	-- 0x1C31
		when 007218 => D <= "11110000";	-- 0x1C32
		when 007219 => D <= "11011001";	-- 0x1C33
		when 007220 => D <= "00100011";	-- 0x1C34
		when 007221 => D <= "11011001";	-- 0x1C35
		when 007222 => D <= "11001001";	-- 0x1C36
		when 007223 => D <= "11101111";	-- 0x1C37
		when 007224 => D <= "11000000";	-- 0x1C38
		when 007225 => D <= "00000010";	-- 0x1C39
		when 007226 => D <= "00101101";	-- 0x1C3A
		when 007227 => D <= "11100000";	-- 0x1C3B
		when 007228 => D <= "00000101";	-- 0x1C3C
		when 007229 => D <= "00100100";	-- 0x1C3D
		when 007230 => D <= "11100000";	-- 0x1C3E
		when 007231 => D <= "00000001";	-- 0x1C3F
		when 007232 => D <= "11000000";	-- 0x1C40
		when 007233 => D <= "00000100";	-- 0x1C41
		when 007234 => D <= "00000011";	-- 0x1C42
		when 007235 => D <= "11100000";	-- 0x1C43
		when 007236 => D <= "00110100";	-- 0x1C44
		when 007237 => D <= "11001001";	-- 0x1C45
		when 007238 => D <= "11101111";	-- 0x1C46
		when 007239 => D <= "00101101";	-- 0x1C47
		when 007240 => D <= "00110010";	-- 0x1C48
		when 007241 => D <= "00000000";	-- 0x1C49
		when 007242 => D <= "00000100";	-- 0x1C4A
		when 007243 => D <= "00110110";	-- 0x1C4B
		when 007244 => D <= "00110100";	-- 0x1C4C
		when 007245 => D <= "11001001";	-- 0x1C4D
		when 007246 => D <= "00101101";	-- 0x1C4E
		when 007247 => D <= "00110110";	-- 0x1C4F
		when 007248 => D <= "11000000";	-- 0x1C50
		when 007249 => D <= "00000011";	-- 0x1C51
		when 007250 => D <= "11100000";	-- 0x1C52
		when 007251 => D <= "00000001";	-- 0x1C53
		when 007252 => D <= "00101100";	-- 0x1C54
		when 007253 => D <= "00000000";	-- 0x1C55
		when 007254 => D <= "00000011";	-- 0x1C56
		when 007255 => D <= "10100001";	-- 0x1C57
		when 007256 => D <= "00000011";	-- 0x1C58
		when 007257 => D <= "00110100";	-- 0x1C59
		when 007258 => D <= "11001001";	-- 0x1C5A
		when 007259 => D <= "11101111";	-- 0x1C5B
		when 007260 => D <= "00110000";	-- 0x1C5C
		when 007261 => D <= "11110001";	-- 0x1C5D
		when 007262 => D <= "00111000";	-- 0x1C5E
		when 007263 => D <= "10101010";	-- 0x1C5F
		when 007264 => D <= "00111011";	-- 0x1C60
		when 007265 => D <= "00101001";	-- 0x1C61
		when 007266 => D <= "00000100";	-- 0x1C62
		when 007267 => D <= "00101101";	-- 0x1C63
		when 007268 => D <= "00100100";	-- 0x1C64
		when 007269 => D <= "11000011";	-- 0x1C65
		when 007270 => D <= "00000011";	-- 0x1C66
		when 007271 => D <= "00101101";	-- 0x1C67
		when 007272 => D <= "00001111";	-- 0x1C68
		when 007273 => D <= "10100001";	-- 0x1C69
		when 007274 => D <= "00000011";	-- 0x1C6A
		when 007275 => D <= "10001000";	-- 0x1C6B
		when 007276 => D <= "00010011";	-- 0x1C6C
		when 007277 => D <= "00110110";	-- 0x1C6D
		when 007278 => D <= "01011000";	-- 0x1C6E
		when 007279 => D <= "01100101";	-- 0x1C6F
		when 007280 => D <= "01100110";	-- 0x1C70
		when 007281 => D <= "10011101";	-- 0x1C71
		when 007282 => D <= "01111000";	-- 0x1C72
		when 007283 => D <= "01100101";	-- 0x1C73
		when 007284 => D <= "01000000";	-- 0x1C74
		when 007285 => D <= "10100010";	-- 0x1C75
		when 007286 => D <= "01100000";	-- 0x1C76
		when 007287 => D <= "00110010";	-- 0x1C77
		when 007288 => D <= "11001001";	-- 0x1C78
		when 007289 => D <= "11100111";	-- 0x1C79
		when 007290 => D <= "00100001";	-- 0x1C7A
		when 007291 => D <= "11110111";	-- 0x1C7B
		when 007292 => D <= "10101111";	-- 0x1C7C
		when 007293 => D <= "00100100";	-- 0x1C7D
		when 007294 => D <= "11101011";	-- 0x1C7E
		when 007295 => D <= "00101111";	-- 0x1C7F
		when 007296 => D <= "10110000";	-- 0x1C80
		when 007297 => D <= "10110000";	-- 0x1C81
		when 007298 => D <= "00010100";	-- 0x1C82
		when 007299 => D <= "11101110";	-- 0x1C83
		when 007300 => D <= "01111110";	-- 0x1C84
		when 007301 => D <= "10111011";	-- 0x1C85
		when 007302 => D <= "10010100";	-- 0x1C86
		when 007303 => D <= "01011000";	-- 0x1C87
		when 007304 => D <= "11110001";	-- 0x1C88
		when 007305 => D <= "00111010";	-- 0x1C89
		when 007306 => D <= "01111110";	-- 0x1C8A
		when 007307 => D <= "11111000";	-- 0x1C8B
		when 007308 => D <= "11001111";	-- 0x1C8C
		when 007309 => D <= "11100011";	-- 0x1C8D
		when 007310 => D <= "00110100";	-- 0x1C8E
		when 007311 => D <= "11001101";	-- 0x1C8F
		when 007312 => D <= "11001101";	-- 0x1C90
		when 007313 => D <= "00010101";	-- 0x1C91
		when 007314 => D <= "00100000";	-- 0x1C92
		when 007315 => D <= "00000111";	-- 0x1C93
		when 007316 => D <= "00111000";	-- 0x1C94
		when 007317 => D <= "00000011";	-- 0x1C95
		when 007318 => D <= "10000110";	-- 0x1C96
		when 007319 => D <= "00110000";	-- 0x1C97
		when 007320 => D <= "00001001";	-- 0x1C98
		when 007321 => D <= "11001111";	-- 0x1C99
		when 007322 => D <= "00000101";	-- 0x1C9A
		when 007323 => D <= "00111000";	-- 0x1C9B
		when 007324 => D <= "00000111";	-- 0x1C9C
		when 007325 => D <= "10010110";	-- 0x1C9D
		when 007326 => D <= "00110000";	-- 0x1C9E
		when 007327 => D <= "00000100";	-- 0x1C9F
		when 007328 => D <= "11101101";	-- 0x1CA0
		when 007329 => D <= "01000100";	-- 0x1CA1
		when 007330 => D <= "01110111";	-- 0x1CA2
		when 007331 => D <= "11001001";	-- 0x1CA3
		when 007332 => D <= "11101111";	-- 0x1CA4
		when 007333 => D <= "00000010";	-- 0x1CA5
		when 007334 => D <= "10100000";	-- 0x1CA6
		when 007335 => D <= "00110100";	-- 0x1CA7
		when 007336 => D <= "11001001";	-- 0x1CA8
		when 007337 => D <= "11101111";	-- 0x1CA9
		when 007338 => D <= "00101101";	-- 0x1CAA
		when 007339 => D <= "00110011";	-- 0x1CAB
		when 007340 => D <= "00000000";	-- 0x1CAC
		when 007341 => D <= "00000100";	-- 0x1CAD
		when 007342 => D <= "00110100";	-- 0x1CAE
		when 007343 => D <= "11001111";	-- 0x1CAF
		when 007344 => D <= "00001001";	-- 0x1CB0
		when 007345 => D <= "10100000";	-- 0x1CB1
		when 007346 => D <= "00000010";	-- 0x1CB2
		when 007347 => D <= "00110100";	-- 0x1CB3
		when 007348 => D <= "01111110";	-- 0x1CB4
		when 007349 => D <= "00110110";	-- 0x1CB5
		when 007350 => D <= "10000000";	-- 0x1CB6
		when 007351 => D <= "11001101";	-- 0x1CB7
		when 007352 => D <= "00011101";	-- 0x1CB8
		when 007353 => D <= "00010101";	-- 0x1CB9
		when 007354 => D <= "11101111";	-- 0x1CBA
		when 007355 => D <= "00110000";	-- 0x1CBB
		when 007356 => D <= "00111000";	-- 0x1CBC
		when 007357 => D <= "00000000";	-- 0x1CBD
		when 007358 => D <= "00000011";	-- 0x1CBE
		when 007359 => D <= "00000001";	-- 0x1CBF
		when 007360 => D <= "00101101";	-- 0x1CC0
		when 007361 => D <= "00110000";	-- 0x1CC1
		when 007362 => D <= "11110000";	-- 0x1CC2
		when 007363 => D <= "01001100";	-- 0x1CC3
		when 007364 => D <= "11001100";	-- 0x1CC4
		when 007365 => D <= "11001100";	-- 0x1CC5
		when 007366 => D <= "11001101";	-- 0x1CC6
		when 007367 => D <= "00000011";	-- 0x1CC7
		when 007368 => D <= "00110011";	-- 0x1CC8
		when 007369 => D <= "00000000";	-- 0x1CC9
		when 007370 => D <= "00001000";	-- 0x1CCA
		when 007371 => D <= "00000001";	-- 0x1CCB
		when 007372 => D <= "10100001";	-- 0x1CCC
		when 007373 => D <= "00000011";	-- 0x1CCD
		when 007374 => D <= "00000001";	-- 0x1CCE
		when 007375 => D <= "00110100";	-- 0x1CCF
		when 007376 => D <= "00110100";	-- 0x1CD0
		when 007377 => D <= "11101111";	-- 0x1CD1
		when 007378 => D <= "00000001";	-- 0x1CD2
		when 007379 => D <= "00110000";	-- 0x1CD3
		when 007380 => D <= "11110000";	-- 0x1CD4
		when 007381 => D <= "00110001";	-- 0x1CD5
		when 007382 => D <= "01110010";	-- 0x1CD6
		when 007383 => D <= "00010111";	-- 0x1CD7
		when 007384 => D <= "11111000";	-- 0x1CD8
		when 007385 => D <= "00000100";	-- 0x1CD9
		when 007386 => D <= "00000001";	-- 0x1CDA
		when 007387 => D <= "10100010";	-- 0x1CDB
		when 007388 => D <= "00000011";	-- 0x1CDC
		when 007389 => D <= "10100010";	-- 0x1CDD
		when 007390 => D <= "00000011";	-- 0x1CDE
		when 007391 => D <= "00101101";	-- 0x1CDF
		when 007392 => D <= "00110000";	-- 0x1CE0
		when 007393 => D <= "00110010";	-- 0x1CE1
		when 007394 => D <= "00100000";	-- 0x1CE2
		when 007395 => D <= "00000100";	-- 0x1CE3
		when 007396 => D <= "10100010";	-- 0x1CE4
		when 007397 => D <= "00000011";	-- 0x1CE5
		when 007398 => D <= "10001100";	-- 0x1CE6
		when 007399 => D <= "00010001";	-- 0x1CE7
		when 007400 => D <= "10101100";	-- 0x1CE8
		when 007401 => D <= "00010100";	-- 0x1CE9
		when 007402 => D <= "00001001";	-- 0x1CEA
		when 007403 => D <= "01010110";	-- 0x1CEB
		when 007404 => D <= "11011010";	-- 0x1CEC
		when 007405 => D <= "10100101";	-- 0x1CED
		when 007406 => D <= "01011001";	-- 0x1CEE
		when 007407 => D <= "00110000";	-- 0x1CEF
		when 007408 => D <= "11000101";	-- 0x1CF0
		when 007409 => D <= "01011100";	-- 0x1CF1
		when 007410 => D <= "10010000";	-- 0x1CF2
		when 007411 => D <= "10101010";	-- 0x1CF3
		when 007412 => D <= "10011110";	-- 0x1CF4
		when 007413 => D <= "01110000";	-- 0x1CF5
		when 007414 => D <= "01101111";	-- 0x1CF6
		when 007415 => D <= "01100001";	-- 0x1CF7
		when 007416 => D <= "10100001";	-- 0x1CF8
		when 007417 => D <= "11001011";	-- 0x1CF9
		when 007418 => D <= "11011010";	-- 0x1CFA
		when 007419 => D <= "10010110";	-- 0x1CFB
		when 007420 => D <= "10100100";	-- 0x1CFC
		when 007421 => D <= "00110001";	-- 0x1CFD
		when 007422 => D <= "10011111";	-- 0x1CFE
		when 007423 => D <= "10110100";	-- 0x1CFF
		when 007424 => D <= "11100111";	-- 0x1D00
		when 007425 => D <= "10100000";	-- 0x1D01
		when 007426 => D <= "11111110";	-- 0x1D02
		when 007427 => D <= "01011100";	-- 0x1D03
		when 007428 => D <= "11111100";	-- 0x1D04
		when 007429 => D <= "11101010";	-- 0x1D05
		when 007430 => D <= "00011011";	-- 0x1D06
		when 007431 => D <= "01000011";	-- 0x1D07
		when 007432 => D <= "11001010";	-- 0x1D08
		when 007433 => D <= "00110110";	-- 0x1D09
		when 007434 => D <= "11101101";	-- 0x1D0A
		when 007435 => D <= "10100111";	-- 0x1D0B
		when 007436 => D <= "10011100";	-- 0x1D0C
		when 007437 => D <= "01111110";	-- 0x1D0D
		when 007438 => D <= "01011110";	-- 0x1D0E
		when 007439 => D <= "11110000";	-- 0x1D0F
		when 007440 => D <= "01101110";	-- 0x1D10
		when 007441 => D <= "00100011";	-- 0x1D11
		when 007442 => D <= "10000000";	-- 0x1D12
		when 007443 => D <= "10010011";	-- 0x1D13
		when 007444 => D <= "00000100";	-- 0x1D14
		when 007445 => D <= "00001111";	-- 0x1D15
		when 007446 => D <= "00110100";	-- 0x1D16
		when 007447 => D <= "11001001";	-- 0x1D17
		when 007448 => D <= "11101111";	-- 0x1D18
		when 007449 => D <= "00110000";	-- 0x1D19
		when 007450 => D <= "11101110";	-- 0x1D1A
		when 007451 => D <= "00100010";	-- 0x1D1B
		when 007452 => D <= "11111001";	-- 0x1D1C
		when 007453 => D <= "10000011";	-- 0x1D1D
		when 007454 => D <= "01101110";	-- 0x1D1E
		when 007455 => D <= "00000100";	-- 0x1D1F
		when 007456 => D <= "00101101";	-- 0x1D20
		when 007457 => D <= "10100010";	-- 0x1D21
		when 007458 => D <= "00001111";	-- 0x1D22
		when 007459 => D <= "00100100";	-- 0x1D23
		when 007460 => D <= "00000011";	-- 0x1D24
		when 007461 => D <= "00101101";	-- 0x1D25
		when 007462 => D <= "00001111";	-- 0x1D26
		when 007463 => D <= "00101101";	-- 0x1D27
		when 007464 => D <= "00001111";	-- 0x1D28
		when 007465 => D <= "00101101";	-- 0x1D29
		when 007466 => D <= "00100111";	-- 0x1D2A
		when 007467 => D <= "10100001";	-- 0x1D2B
		when 007468 => D <= "00000011";	-- 0x1D2C
		when 007469 => D <= "00101101";	-- 0x1D2D
		when 007470 => D <= "00110011";	-- 0x1D2E
		when 007471 => D <= "11000000";	-- 0x1D2F
		when 007472 => D <= "00000000";	-- 0x1D30
		when 007473 => D <= "00000100";	-- 0x1D31
		when 007474 => D <= "00000010";	-- 0x1D32
		when 007475 => D <= "00110100";	-- 0x1D33
		when 007476 => D <= "11001001";	-- 0x1D34
		when 007477 => D <= "10100001";	-- 0x1D35
		when 007478 => D <= "00000011";	-- 0x1D36
		when 007479 => D <= "00000001";	-- 0x1D37
		when 007480 => D <= "00110010";	-- 0x1D38
		when 007481 => D <= "00000000";	-- 0x1D39
		when 007482 => D <= "00000010";	-- 0x1D3A
		when 007483 => D <= "00011000";	-- 0x1D3B
		when 007484 => D <= "00110100";	-- 0x1D3C
		when 007485 => D <= "11001001";	-- 0x1D3D
		when 007486 => D <= "11101111";	-- 0x1D3E
		when 007487 => D <= "00110101";	-- 0x1D3F
		when 007488 => D <= "00100111";	-- 0x1D40
		when 007489 => D <= "10100001";	-- 0x1D41
		when 007490 => D <= "00000011";	-- 0x1D42
		when 007491 => D <= "11100000";	-- 0x1D43
		when 007492 => D <= "00000000";	-- 0x1D44
		when 007493 => D <= "00000110";	-- 0x1D45
		when 007494 => D <= "00011000";	-- 0x1D46
		when 007495 => D <= "00101111";	-- 0x1D47
		when 007496 => D <= "00000011";	-- 0x1D48
		when 007497 => D <= "11101111";	-- 0x1D49
		when 007498 => D <= "00110101";	-- 0x1D4A
		when 007499 => D <= "00101101";	-- 0x1D4B
		when 007500 => D <= "00101101";	-- 0x1D4C
		when 007501 => D <= "00000100";	-- 0x1D4D
		when 007502 => D <= "00101101";	-- 0x1D4E
		when 007503 => D <= "00001111";	-- 0x1D4F
		when 007504 => D <= "10100001";	-- 0x1D50
		when 007505 => D <= "00000011";	-- 0x1D51
		when 007506 => D <= "10000110";	-- 0x1D52
		when 007507 => D <= "00010100";	-- 0x1D53
		when 007508 => D <= "11100110";	-- 0x1D54
		when 007509 => D <= "01011100";	-- 0x1D55
		when 007510 => D <= "00011111";	-- 0x1D56
		when 007511 => D <= "00001011";	-- 0x1D57
		when 007512 => D <= "10100011";	-- 0x1D58
		when 007513 => D <= "10001111";	-- 0x1D59
		when 007514 => D <= "00111000";	-- 0x1D5A
		when 007515 => D <= "11101110";	-- 0x1D5B
		when 007516 => D <= "11101001";	-- 0x1D5C
		when 007517 => D <= "00010101";	-- 0x1D5D
		when 007518 => D <= "01100011";	-- 0x1D5E
		when 007519 => D <= "10111011";	-- 0x1D5F
		when 007520 => D <= "00100011";	-- 0x1D60
		when 007521 => D <= "11101110";	-- 0x1D61
		when 007522 => D <= "10010010";	-- 0x1D62
		when 007523 => D <= "00001101";	-- 0x1D63
		when 007524 => D <= "11001101";	-- 0x1D64
		when 007525 => D <= "11101101";	-- 0x1D65
		when 007526 => D <= "11110001";	-- 0x1D66
		when 007527 => D <= "00100011";	-- 0x1D67
		when 007528 => D <= "01011101";	-- 0x1D68
		when 007529 => D <= "00011011";	-- 0x1D69
		when 007530 => D <= "11101010";	-- 0x1D6A
		when 007531 => D <= "00000100";	-- 0x1D6B
		when 007532 => D <= "00110100";	-- 0x1D6C
		when 007533 => D <= "11001001";	-- 0x1D6D
		when 007534 => D <= "11101111";	-- 0x1D6E
		when 007535 => D <= "00101101";	-- 0x1D6F
		when 007536 => D <= "00011100";	-- 0x1D70
		when 007537 => D <= "00000001";	-- 0x1D71
		when 007538 => D <= "00011101";	-- 0x1D72
		when 007539 => D <= "00000101";	-- 0x1D73
		when 007540 => D <= "00110100";	-- 0x1D74
		when 007541 => D <= "11001001";	-- 0x1D75
		when 007542 => D <= "01111110";	-- 0x1D76
		when 007543 => D <= "11111110";	-- 0x1D77
		when 007544 => D <= "10000001";	-- 0x1D78
		when 007545 => D <= "00111000";	-- 0x1D79
		when 007546 => D <= "00001110";	-- 0x1D7A
		when 007547 => D <= "11101111";	-- 0x1D7B
		when 007548 => D <= "10100001";	-- 0x1D7C
		when 007549 => D <= "00011000";	-- 0x1D7D
		when 007550 => D <= "00000001";	-- 0x1D7E
		when 007551 => D <= "00000101";	-- 0x1D7F
		when 007552 => D <= "00101101";	-- 0x1D80
		when 007553 => D <= "00110010";	-- 0x1D81
		when 007554 => D <= "10100011";	-- 0x1D82
		when 007555 => D <= "00000001";	-- 0x1D83
		when 007556 => D <= "00000000";	-- 0x1D84
		when 007557 => D <= "00000110";	-- 0x1D85
		when 007558 => D <= "00011000";	-- 0x1D86
		when 007559 => D <= "00101111";	-- 0x1D87
		when 007560 => D <= "00000011";	-- 0x1D88
		when 007561 => D <= "11101111";	-- 0x1D89
		when 007562 => D <= "10100000";	-- 0x1D8A
		when 007563 => D <= "00000001";	-- 0x1D8B
		when 007564 => D <= "00101101";	-- 0x1D8C
		when 007565 => D <= "00101101";	-- 0x1D8D
		when 007566 => D <= "00000100";	-- 0x1D8E
		when 007567 => D <= "00101101";	-- 0x1D8F
		when 007568 => D <= "00001111";	-- 0x1D90
		when 007569 => D <= "10100001";	-- 0x1D91
		when 007570 => D <= "00000011";	-- 0x1D92
		when 007571 => D <= "10001100";	-- 0x1D93
		when 007572 => D <= "00010000";	-- 0x1D94
		when 007573 => D <= "10110010";	-- 0x1D95
		when 007574 => D <= "00010011";	-- 0x1D96
		when 007575 => D <= "00001110";	-- 0x1D97
		when 007576 => D <= "01010101";	-- 0x1D98
		when 007577 => D <= "11100100";	-- 0x1D99
		when 007578 => D <= "10001101";	-- 0x1D9A
		when 007579 => D <= "01011000";	-- 0x1D9B
		when 007580 => D <= "00111001";	-- 0x1D9C
		when 007581 => D <= "10111100";	-- 0x1D9D
		when 007582 => D <= "01011011";	-- 0x1D9E
		when 007583 => D <= "10011000";	-- 0x1D9F
		when 007584 => D <= "11111101";	-- 0x1DA0
		when 007585 => D <= "10011110";	-- 0x1DA1
		when 007586 => D <= "00000000";	-- 0x1DA2
		when 007587 => D <= "00110110";	-- 0x1DA3
		when 007588 => D <= "01110101";	-- 0x1DA4
		when 007589 => D <= "10100000";	-- 0x1DA5
		when 007590 => D <= "11011011";	-- 0x1DA6
		when 007591 => D <= "11101000";	-- 0x1DA7
		when 007592 => D <= "10110100";	-- 0x1DA8
		when 007593 => D <= "01100011";	-- 0x1DA9
		when 007594 => D <= "01000010";	-- 0x1DAA
		when 007595 => D <= "11000100";	-- 0x1DAB
		when 007596 => D <= "11100110";	-- 0x1DAC
		when 007597 => D <= "10110101";	-- 0x1DAD
		when 007598 => D <= "00001001";	-- 0x1DAE
		when 007599 => D <= "00110110";	-- 0x1DAF
		when 007600 => D <= "10111110";	-- 0x1DB0
		when 007601 => D <= "11101001";	-- 0x1DB1
		when 007602 => D <= "00110110";	-- 0x1DB2
		when 007603 => D <= "01110011";	-- 0x1DB3
		when 007604 => D <= "00011011";	-- 0x1DB4
		when 007605 => D <= "01011101";	-- 0x1DB5
		when 007606 => D <= "11101100";	-- 0x1DB6
		when 007607 => D <= "11011000";	-- 0x1DB7
		when 007608 => D <= "11011110";	-- 0x1DB8
		when 007609 => D <= "01100011";	-- 0x1DB9
		when 007610 => D <= "10111110";	-- 0x1DBA
		when 007611 => D <= "11110000";	-- 0x1DBB
		when 007612 => D <= "01100001";	-- 0x1DBC
		when 007613 => D <= "10100001";	-- 0x1DBD
		when 007614 => D <= "10110011";	-- 0x1DBE
		when 007615 => D <= "00001100";	-- 0x1DBF
		when 007616 => D <= "00000100";	-- 0x1DC0
		when 007617 => D <= "00001111";	-- 0x1DC1
		when 007618 => D <= "00110100";	-- 0x1DC2
		when 007619 => D <= "11001001";	-- 0x1DC3
		when 007620 => D <= "11101111";	-- 0x1DC4
		when 007621 => D <= "00101101";	-- 0x1DC5
		when 007622 => D <= "00101101";	-- 0x1DC6
		when 007623 => D <= "00000100";	-- 0x1DC7
		when 007624 => D <= "10100001";	-- 0x1DC8
		when 007625 => D <= "00000011";	-- 0x1DC9
		when 007626 => D <= "00011000";	-- 0x1DCA
		when 007627 => D <= "00100101";	-- 0x1DCB
		when 007628 => D <= "10100001";	-- 0x1DCC
		when 007629 => D <= "00001111";	-- 0x1DCD
		when 007630 => D <= "00000101";	-- 0x1DCE
		when 007631 => D <= "00100001";	-- 0x1DCF
		when 007632 => D <= "00101101";	-- 0x1DD0
		when 007633 => D <= "00001111";	-- 0x1DD1
		when 007634 => D <= "00110100";	-- 0x1DD2
		when 007635 => D <= "11001001";	-- 0x1DD3
		when 007636 => D <= "11101111";	-- 0x1DD4
		when 007637 => D <= "00011111";	-- 0x1DD5
		when 007638 => D <= "10100011";	-- 0x1DD6
		when 007639 => D <= "00000011";	-- 0x1DD7
		when 007640 => D <= "00011000";	-- 0x1DD8
		when 007641 => D <= "00110100";	-- 0x1DD9
		when 007642 => D <= "11001001";	-- 0x1DDA
		when 007643 => D <= "11101111";	-- 0x1DDB
		when 007644 => D <= "00101101";	-- 0x1DDC
		when 007645 => D <= "00101100";	-- 0x1DDD
		when 007646 => D <= "00000000";	-- 0x1DDE
		when 007647 => D <= "00011110";	-- 0x1DDF
		when 007648 => D <= "10100010";	-- 0x1DE0
		when 007649 => D <= "00110100";	-- 0x1DE1
		when 007650 => D <= "11101111";	-- 0x1DE2
		when 007651 => D <= "00000001";	-- 0x1DE3
		when 007652 => D <= "00101101";	-- 0x1DE4
		when 007653 => D <= "00101100";	-- 0x1DE5
		when 007654 => D <= "00000000";	-- 0x1DE6
		when 007655 => D <= "00000111";	-- 0x1DE7
		when 007656 => D <= "00100010";	-- 0x1DE8
		when 007657 => D <= "00000100";	-- 0x1DE9
		when 007658 => D <= "00110100";	-- 0x1DEA
		when 007659 => D <= "11000011";	-- 0x1DEB
		when 007660 => D <= "01011011";	-- 0x1DEC
		when 007661 => D <= "00011100";	-- 0x1DED
		when 007662 => D <= "00000010";	-- 0x1DEE
		when 007663 => D <= "00101101";	-- 0x1DEF
		when 007664 => D <= "00101100";	-- 0x1DF0
		when 007665 => D <= "00000000";	-- 0x1DF1
		when 007666 => D <= "00001001";	-- 0x1DF2
		when 007667 => D <= "10100000";	-- 0x1DF3
		when 007668 => D <= "00000001";	-- 0x1DF4
		when 007669 => D <= "00110011";	-- 0x1DF5
		when 007670 => D <= "00000000";	-- 0x1DF6
		when 007671 => D <= "00000110";	-- 0x1DF7
		when 007672 => D <= "10100001";	-- 0x1DF8
		when 007673 => D <= "00000001";	-- 0x1DF9
		when 007674 => D <= "00000101";	-- 0x1DFA
		when 007675 => D <= "00000010";	-- 0x1DFB
		when 007676 => D <= "10100001";	-- 0x1DFC
		when 007677 => D <= "00110100";	-- 0x1DFD
		when 007678 => D <= "11001001";	-- 0x1DFE
		when 007679 => D <= "11111111";	-- 0x1DFF
		when 007680 => D <= "00000000";	-- 0x1E00
		when 007681 => D <= "00000000";	-- 0x1E01
		when 007682 => D <= "00000000";	-- 0x1E02
		when 007683 => D <= "00000000";	-- 0x1E03
		when 007684 => D <= "00000000";	-- 0x1E04
		when 007685 => D <= "00000000";	-- 0x1E05
		when 007686 => D <= "00000000";	-- 0x1E06
		when 007687 => D <= "00000000";	-- 0x1E07
		when 007688 => D <= "11110000";	-- 0x1E08
		when 007689 => D <= "11110000";	-- 0x1E09
		when 007690 => D <= "11110000";	-- 0x1E0A
		when 007691 => D <= "11110000";	-- 0x1E0B
		when 007692 => D <= "00000000";	-- 0x1E0C
		when 007693 => D <= "00000000";	-- 0x1E0D
		when 007694 => D <= "00000000";	-- 0x1E0E
		when 007695 => D <= "00000000";	-- 0x1E0F
		when 007696 => D <= "00001111";	-- 0x1E10
		when 007697 => D <= "00001111";	-- 0x1E11
		when 007698 => D <= "00001111";	-- 0x1E12
		when 007699 => D <= "00001111";	-- 0x1E13
		when 007700 => D <= "00000000";	-- 0x1E14
		when 007701 => D <= "00000000";	-- 0x1E15
		when 007702 => D <= "00000000";	-- 0x1E16
		when 007703 => D <= "00000000";	-- 0x1E17
		when 007704 => D <= "11111111";	-- 0x1E18
		when 007705 => D <= "11111111";	-- 0x1E19
		when 007706 => D <= "11111111";	-- 0x1E1A
		when 007707 => D <= "11111111";	-- 0x1E1B
		when 007708 => D <= "00000000";	-- 0x1E1C
		when 007709 => D <= "00000000";	-- 0x1E1D
		when 007710 => D <= "00000000";	-- 0x1E1E
		when 007711 => D <= "00000000";	-- 0x1E1F
		when 007712 => D <= "00000000";	-- 0x1E20
		when 007713 => D <= "00000000";	-- 0x1E21
		when 007714 => D <= "00000000";	-- 0x1E22
		when 007715 => D <= "00000000";	-- 0x1E23
		when 007716 => D <= "11110000";	-- 0x1E24
		when 007717 => D <= "11110000";	-- 0x1E25
		when 007718 => D <= "11110000";	-- 0x1E26
		when 007719 => D <= "11110000";	-- 0x1E27
		when 007720 => D <= "11110000";	-- 0x1E28
		when 007721 => D <= "11110000";	-- 0x1E29
		when 007722 => D <= "11110000";	-- 0x1E2A
		when 007723 => D <= "11110000";	-- 0x1E2B
		when 007724 => D <= "11110000";	-- 0x1E2C
		when 007725 => D <= "11110000";	-- 0x1E2D
		when 007726 => D <= "11110000";	-- 0x1E2E
		when 007727 => D <= "11110000";	-- 0x1E2F
		when 007728 => D <= "00001111";	-- 0x1E30
		when 007729 => D <= "00001111";	-- 0x1E31
		when 007730 => D <= "00001111";	-- 0x1E32
		when 007731 => D <= "00001111";	-- 0x1E33
		when 007732 => D <= "11110000";	-- 0x1E34
		when 007733 => D <= "11110000";	-- 0x1E35
		when 007734 => D <= "11110000";	-- 0x1E36
		when 007735 => D <= "11110000";	-- 0x1E37
		when 007736 => D <= "11111111";	-- 0x1E38
		when 007737 => D <= "11111111";	-- 0x1E39
		when 007738 => D <= "11111111";	-- 0x1E3A
		when 007739 => D <= "11111111";	-- 0x1E3B
		when 007740 => D <= "11110000";	-- 0x1E3C
		when 007741 => D <= "11110000";	-- 0x1E3D
		when 007742 => D <= "11110000";	-- 0x1E3E
		when 007743 => D <= "11110000";	-- 0x1E3F
		when 007744 => D <= "10101010";	-- 0x1E40
		when 007745 => D <= "01010101";	-- 0x1E41
		when 007746 => D <= "10101010";	-- 0x1E42
		when 007747 => D <= "01010101";	-- 0x1E43
		when 007748 => D <= "10101010";	-- 0x1E44
		when 007749 => D <= "01010101";	-- 0x1E45
		when 007750 => D <= "10101010";	-- 0x1E46
		when 007751 => D <= "01010101";	-- 0x1E47
		when 007752 => D <= "00000000";	-- 0x1E48
		when 007753 => D <= "00000000";	-- 0x1E49
		when 007754 => D <= "00000000";	-- 0x1E4A
		when 007755 => D <= "00000000";	-- 0x1E4B
		when 007756 => D <= "10101010";	-- 0x1E4C
		when 007757 => D <= "01010101";	-- 0x1E4D
		when 007758 => D <= "10101010";	-- 0x1E4E
		when 007759 => D <= "01010101";	-- 0x1E4F
		when 007760 => D <= "10101010";	-- 0x1E50
		when 007761 => D <= "01010101";	-- 0x1E51
		when 007762 => D <= "10101010";	-- 0x1E52
		when 007763 => D <= "01010101";	-- 0x1E53
		when 007764 => D <= "00000000";	-- 0x1E54
		when 007765 => D <= "00000000";	-- 0x1E55
		when 007766 => D <= "00000000";	-- 0x1E56
		when 007767 => D <= "00000000";	-- 0x1E57
		when 007768 => D <= "00000000";	-- 0x1E58
		when 007769 => D <= "00100100";	-- 0x1E59
		when 007770 => D <= "00100100";	-- 0x1E5A
		when 007771 => D <= "00000000";	-- 0x1E5B
		when 007772 => D <= "00000000";	-- 0x1E5C
		when 007773 => D <= "00000000";	-- 0x1E5D
		when 007774 => D <= "00000000";	-- 0x1E5E
		when 007775 => D <= "00000000";	-- 0x1E5F
		when 007776 => D <= "00000000";	-- 0x1E60
		when 007777 => D <= "00011100";	-- 0x1E61
		when 007778 => D <= "00100010";	-- 0x1E62
		when 007779 => D <= "01111000";	-- 0x1E63
		when 007780 => D <= "00100000";	-- 0x1E64
		when 007781 => D <= "00100000";	-- 0x1E65
		when 007782 => D <= "01111110";	-- 0x1E66
		when 007783 => D <= "00000000";	-- 0x1E67
		when 007784 => D <= "00000000";	-- 0x1E68
		when 007785 => D <= "00001000";	-- 0x1E69
		when 007786 => D <= "00111110";	-- 0x1E6A
		when 007787 => D <= "00101000";	-- 0x1E6B
		when 007788 => D <= "00111110";	-- 0x1E6C
		when 007789 => D <= "00001010";	-- 0x1E6D
		when 007790 => D <= "00111110";	-- 0x1E6E
		when 007791 => D <= "00001000";	-- 0x1E6F
		when 007792 => D <= "00000000";	-- 0x1E70
		when 007793 => D <= "00000000";	-- 0x1E71
		when 007794 => D <= "00000000";	-- 0x1E72
		when 007795 => D <= "00010000";	-- 0x1E73
		when 007796 => D <= "00000000";	-- 0x1E74
		when 007797 => D <= "00000000";	-- 0x1E75
		when 007798 => D <= "00010000";	-- 0x1E76
		when 007799 => D <= "00000000";	-- 0x1E77
		when 007800 => D <= "00000000";	-- 0x1E78
		when 007801 => D <= "00111100";	-- 0x1E79
		when 007802 => D <= "01000010";	-- 0x1E7A
		when 007803 => D <= "00000100";	-- 0x1E7B
		when 007804 => D <= "00001000";	-- 0x1E7C
		when 007805 => D <= "00000000";	-- 0x1E7D
		when 007806 => D <= "00001000";	-- 0x1E7E
		when 007807 => D <= "00000000";	-- 0x1E7F
		when 007808 => D <= "00000000";	-- 0x1E80
		when 007809 => D <= "00000100";	-- 0x1E81
		when 007810 => D <= "00001000";	-- 0x1E82
		when 007811 => D <= "00001000";	-- 0x1E83
		when 007812 => D <= "00001000";	-- 0x1E84
		when 007813 => D <= "00001000";	-- 0x1E85
		when 007814 => D <= "00000100";	-- 0x1E86
		when 007815 => D <= "00000000";	-- 0x1E87
		when 007816 => D <= "00000000";	-- 0x1E88
		when 007817 => D <= "00100000";	-- 0x1E89
		when 007818 => D <= "00010000";	-- 0x1E8A
		when 007819 => D <= "00010000";	-- 0x1E8B
		when 007820 => D <= "00010000";	-- 0x1E8C
		when 007821 => D <= "00010000";	-- 0x1E8D
		when 007822 => D <= "00100000";	-- 0x1E8E
		when 007823 => D <= "00000000";	-- 0x1E8F
		when 007824 => D <= "00000000";	-- 0x1E90
		when 007825 => D <= "00000000";	-- 0x1E91
		when 007826 => D <= "00010000";	-- 0x1E92
		when 007827 => D <= "00001000";	-- 0x1E93
		when 007828 => D <= "00000100";	-- 0x1E94
		when 007829 => D <= "00001000";	-- 0x1E95
		when 007830 => D <= "00010000";	-- 0x1E96
		when 007831 => D <= "00000000";	-- 0x1E97
		when 007832 => D <= "00000000";	-- 0x1E98
		when 007833 => D <= "00000000";	-- 0x1E99
		when 007834 => D <= "00000100";	-- 0x1E9A
		when 007835 => D <= "00001000";	-- 0x1E9B
		when 007836 => D <= "00010000";	-- 0x1E9C
		when 007837 => D <= "00001000";	-- 0x1E9D
		when 007838 => D <= "00000100";	-- 0x1E9E
		when 007839 => D <= "00000000";	-- 0x1E9F
		when 007840 => D <= "00000000";	-- 0x1EA0
		when 007841 => D <= "00000000";	-- 0x1EA1
		when 007842 => D <= "00000000";	-- 0x1EA2
		when 007843 => D <= "00111110";	-- 0x1EA3
		when 007844 => D <= "00000000";	-- 0x1EA4
		when 007845 => D <= "00111110";	-- 0x1EA5
		when 007846 => D <= "00000000";	-- 0x1EA6
		when 007847 => D <= "00000000";	-- 0x1EA7
		when 007848 => D <= "00000000";	-- 0x1EA8
		when 007849 => D <= "00000000";	-- 0x1EA9
		when 007850 => D <= "00001000";	-- 0x1EAA
		when 007851 => D <= "00001000";	-- 0x1EAB
		when 007852 => D <= "00111110";	-- 0x1EAC
		when 007853 => D <= "00001000";	-- 0x1EAD
		when 007854 => D <= "00001000";	-- 0x1EAE
		when 007855 => D <= "00000000";	-- 0x1EAF
		when 007856 => D <= "00000000";	-- 0x1EB0
		when 007857 => D <= "00000000";	-- 0x1EB1
		when 007858 => D <= "00000000";	-- 0x1EB2
		when 007859 => D <= "00000000";	-- 0x1EB3
		when 007860 => D <= "00111110";	-- 0x1EB4
		when 007861 => D <= "00000000";	-- 0x1EB5
		when 007862 => D <= "00000000";	-- 0x1EB6
		when 007863 => D <= "00000000";	-- 0x1EB7
		when 007864 => D <= "00000000";	-- 0x1EB8
		when 007865 => D <= "00000000";	-- 0x1EB9
		when 007866 => D <= "00010100";	-- 0x1EBA
		when 007867 => D <= "00001000";	-- 0x1EBB
		when 007868 => D <= "00111110";	-- 0x1EBC
		when 007869 => D <= "00001000";	-- 0x1EBD
		when 007870 => D <= "00010100";	-- 0x1EBE
		when 007871 => D <= "00000000";	-- 0x1EBF
		when 007872 => D <= "00000000";	-- 0x1EC0
		when 007873 => D <= "00000000";	-- 0x1EC1
		when 007874 => D <= "00000010";	-- 0x1EC2
		when 007875 => D <= "00000100";	-- 0x1EC3
		when 007876 => D <= "00001000";	-- 0x1EC4
		when 007877 => D <= "00010000";	-- 0x1EC5
		when 007878 => D <= "00100000";	-- 0x1EC6
		when 007879 => D <= "00000000";	-- 0x1EC7
		when 007880 => D <= "00000000";	-- 0x1EC8
		when 007881 => D <= "00000000";	-- 0x1EC9
		when 007882 => D <= "00010000";	-- 0x1ECA
		when 007883 => D <= "00000000";	-- 0x1ECB
		when 007884 => D <= "00000000";	-- 0x1ECC
		when 007885 => D <= "00010000";	-- 0x1ECD
		when 007886 => D <= "00010000";	-- 0x1ECE
		when 007887 => D <= "00100000";	-- 0x1ECF
		when 007888 => D <= "00000000";	-- 0x1ED0
		when 007889 => D <= "00000000";	-- 0x1ED1
		when 007890 => D <= "00000000";	-- 0x1ED2
		when 007891 => D <= "00000000";	-- 0x1ED3
		when 007892 => D <= "00000000";	-- 0x1ED4
		when 007893 => D <= "00001000";	-- 0x1ED5
		when 007894 => D <= "00001000";	-- 0x1ED6
		when 007895 => D <= "00010000";	-- 0x1ED7
		when 007896 => D <= "00000000";	-- 0x1ED8
		when 007897 => D <= "00000000";	-- 0x1ED9
		when 007898 => D <= "00000000";	-- 0x1EDA
		when 007899 => D <= "00000000";	-- 0x1EDB
		when 007900 => D <= "00000000";	-- 0x1EDC
		when 007901 => D <= "00011000";	-- 0x1EDD
		when 007902 => D <= "00011000";	-- 0x1EDE
		when 007903 => D <= "00000000";	-- 0x1EDF
		when 007904 => D <= "00000000";	-- 0x1EE0
		when 007905 => D <= "00111100";	-- 0x1EE1
		when 007906 => D <= "01000110";	-- 0x1EE2
		when 007907 => D <= "01001010";	-- 0x1EE3
		when 007908 => D <= "01010010";	-- 0x1EE4
		when 007909 => D <= "01100010";	-- 0x1EE5
		when 007910 => D <= "00111100";	-- 0x1EE6
		when 007911 => D <= "00000000";	-- 0x1EE7
		when 007912 => D <= "00000000";	-- 0x1EE8
		when 007913 => D <= "00011000";	-- 0x1EE9
		when 007914 => D <= "00101000";	-- 0x1EEA
		when 007915 => D <= "00001000";	-- 0x1EEB
		when 007916 => D <= "00001000";	-- 0x1EEC
		when 007917 => D <= "00001000";	-- 0x1EED
		when 007918 => D <= "00111110";	-- 0x1EEE
		when 007919 => D <= "00000000";	-- 0x1EEF
		when 007920 => D <= "00000000";	-- 0x1EF0
		when 007921 => D <= "00111100";	-- 0x1EF1
		when 007922 => D <= "01000010";	-- 0x1EF2
		when 007923 => D <= "00000010";	-- 0x1EF3
		when 007924 => D <= "00111100";	-- 0x1EF4
		when 007925 => D <= "01000000";	-- 0x1EF5
		when 007926 => D <= "01111110";	-- 0x1EF6
		when 007927 => D <= "00000000";	-- 0x1EF7
		when 007928 => D <= "00000000";	-- 0x1EF8
		when 007929 => D <= "00111100";	-- 0x1EF9
		when 007930 => D <= "01000010";	-- 0x1EFA
		when 007931 => D <= "00001100";	-- 0x1EFB
		when 007932 => D <= "00000010";	-- 0x1EFC
		when 007933 => D <= "01000010";	-- 0x1EFD
		when 007934 => D <= "00111100";	-- 0x1EFE
		when 007935 => D <= "00000000";	-- 0x1EFF
		when 007936 => D <= "00000000";	-- 0x1F00
		when 007937 => D <= "00001000";	-- 0x1F01
		when 007938 => D <= "00011000";	-- 0x1F02
		when 007939 => D <= "00101000";	-- 0x1F03
		when 007940 => D <= "01001000";	-- 0x1F04
		when 007941 => D <= "01111110";	-- 0x1F05
		when 007942 => D <= "00001000";	-- 0x1F06
		when 007943 => D <= "00000000";	-- 0x1F07
		when 007944 => D <= "00000000";	-- 0x1F08
		when 007945 => D <= "01111110";	-- 0x1F09
		when 007946 => D <= "01000000";	-- 0x1F0A
		when 007947 => D <= "01111100";	-- 0x1F0B
		when 007948 => D <= "00000010";	-- 0x1F0C
		when 007949 => D <= "01000010";	-- 0x1F0D
		when 007950 => D <= "00111100";	-- 0x1F0E
		when 007951 => D <= "00000000";	-- 0x1F0F
		when 007952 => D <= "00000000";	-- 0x1F10
		when 007953 => D <= "00111100";	-- 0x1F11
		when 007954 => D <= "01000000";	-- 0x1F12
		when 007955 => D <= "01111100";	-- 0x1F13
		when 007956 => D <= "01000010";	-- 0x1F14
		when 007957 => D <= "01000010";	-- 0x1F15
		when 007958 => D <= "00111100";	-- 0x1F16
		when 007959 => D <= "00000000";	-- 0x1F17
		when 007960 => D <= "00000000";	-- 0x1F18
		when 007961 => D <= "01111110";	-- 0x1F19
		when 007962 => D <= "00000010";	-- 0x1F1A
		when 007963 => D <= "00000100";	-- 0x1F1B
		when 007964 => D <= "00001000";	-- 0x1F1C
		when 007965 => D <= "00010000";	-- 0x1F1D
		when 007966 => D <= "00010000";	-- 0x1F1E
		when 007967 => D <= "00000000";	-- 0x1F1F
		when 007968 => D <= "00000000";	-- 0x1F20
		when 007969 => D <= "00111100";	-- 0x1F21
		when 007970 => D <= "01000010";	-- 0x1F22
		when 007971 => D <= "00111100";	-- 0x1F23
		when 007972 => D <= "01000010";	-- 0x1F24
		when 007973 => D <= "01000010";	-- 0x1F25
		when 007974 => D <= "00111100";	-- 0x1F26
		when 007975 => D <= "00000000";	-- 0x1F27
		when 007976 => D <= "00000000";	-- 0x1F28
		when 007977 => D <= "00111100";	-- 0x1F29
		when 007978 => D <= "01000010";	-- 0x1F2A
		when 007979 => D <= "01000010";	-- 0x1F2B
		when 007980 => D <= "00111110";	-- 0x1F2C
		when 007981 => D <= "00000010";	-- 0x1F2D
		when 007982 => D <= "00111100";	-- 0x1F2E
		when 007983 => D <= "00000000";	-- 0x1F2F
		when 007984 => D <= "00000000";	-- 0x1F30
		when 007985 => D <= "00111100";	-- 0x1F31
		when 007986 => D <= "01000010";	-- 0x1F32
		when 007987 => D <= "01000010";	-- 0x1F33
		when 007988 => D <= "01111110";	-- 0x1F34
		when 007989 => D <= "01000010";	-- 0x1F35
		when 007990 => D <= "01000010";	-- 0x1F36
		when 007991 => D <= "00000000";	-- 0x1F37
		when 007992 => D <= "00000000";	-- 0x1F38
		when 007993 => D <= "01111100";	-- 0x1F39
		when 007994 => D <= "01000010";	-- 0x1F3A
		when 007995 => D <= "01111100";	-- 0x1F3B
		when 007996 => D <= "01000010";	-- 0x1F3C
		when 007997 => D <= "01000010";	-- 0x1F3D
		when 007998 => D <= "01111100";	-- 0x1F3E
		when 007999 => D <= "00000000";	-- 0x1F3F
		when 008000 => D <= "00000000";	-- 0x1F40
		when 008001 => D <= "00111100";	-- 0x1F41
		when 008002 => D <= "01000010";	-- 0x1F42
		when 008003 => D <= "01000000";	-- 0x1F43
		when 008004 => D <= "01000000";	-- 0x1F44
		when 008005 => D <= "01000010";	-- 0x1F45
		when 008006 => D <= "00111100";	-- 0x1F46
		when 008007 => D <= "00000000";	-- 0x1F47
		when 008008 => D <= "00000000";	-- 0x1F48
		when 008009 => D <= "01111000";	-- 0x1F49
		when 008010 => D <= "01000100";	-- 0x1F4A
		when 008011 => D <= "01000010";	-- 0x1F4B
		when 008012 => D <= "01000010";	-- 0x1F4C
		when 008013 => D <= "01000100";	-- 0x1F4D
		when 008014 => D <= "01111000";	-- 0x1F4E
		when 008015 => D <= "00000000";	-- 0x1F4F
		when 008016 => D <= "00000000";	-- 0x1F50
		when 008017 => D <= "01111110";	-- 0x1F51
		when 008018 => D <= "01000000";	-- 0x1F52
		when 008019 => D <= "01111100";	-- 0x1F53
		when 008020 => D <= "01000000";	-- 0x1F54
		when 008021 => D <= "01000000";	-- 0x1F55
		when 008022 => D <= "01111110";	-- 0x1F56
		when 008023 => D <= "00000000";	-- 0x1F57
		when 008024 => D <= "00000000";	-- 0x1F58
		when 008025 => D <= "01111110";	-- 0x1F59
		when 008026 => D <= "01000000";	-- 0x1F5A
		when 008027 => D <= "01111100";	-- 0x1F5B
		when 008028 => D <= "01000000";	-- 0x1F5C
		when 008029 => D <= "01000000";	-- 0x1F5D
		when 008030 => D <= "01000000";	-- 0x1F5E
		when 008031 => D <= "00000000";	-- 0x1F5F
		when 008032 => D <= "00000000";	-- 0x1F60
		when 008033 => D <= "00111100";	-- 0x1F61
		when 008034 => D <= "01000010";	-- 0x1F62
		when 008035 => D <= "01000000";	-- 0x1F63
		when 008036 => D <= "01001110";	-- 0x1F64
		when 008037 => D <= "01000010";	-- 0x1F65
		when 008038 => D <= "00111100";	-- 0x1F66
		when 008039 => D <= "00000000";	-- 0x1F67
		when 008040 => D <= "00000000";	-- 0x1F68
		when 008041 => D <= "01000010";	-- 0x1F69
		when 008042 => D <= "01000010";	-- 0x1F6A
		when 008043 => D <= "01111110";	-- 0x1F6B
		when 008044 => D <= "01000010";	-- 0x1F6C
		when 008045 => D <= "01000010";	-- 0x1F6D
		when 008046 => D <= "01000010";	-- 0x1F6E
		when 008047 => D <= "00000000";	-- 0x1F6F
		when 008048 => D <= "00000000";	-- 0x1F70
		when 008049 => D <= "00111110";	-- 0x1F71
		when 008050 => D <= "00001000";	-- 0x1F72
		when 008051 => D <= "00001000";	-- 0x1F73
		when 008052 => D <= "00001000";	-- 0x1F74
		when 008053 => D <= "00001000";	-- 0x1F75
		when 008054 => D <= "00111110";	-- 0x1F76
		when 008055 => D <= "00000000";	-- 0x1F77
		when 008056 => D <= "00000000";	-- 0x1F78
		when 008057 => D <= "00000010";	-- 0x1F79
		when 008058 => D <= "00000010";	-- 0x1F7A
		when 008059 => D <= "00000010";	-- 0x1F7B
		when 008060 => D <= "01000010";	-- 0x1F7C
		when 008061 => D <= "01000010";	-- 0x1F7D
		when 008062 => D <= "00111100";	-- 0x1F7E
		when 008063 => D <= "00000000";	-- 0x1F7F
		when 008064 => D <= "00000000";	-- 0x1F80
		when 008065 => D <= "01000100";	-- 0x1F81
		when 008066 => D <= "01001000";	-- 0x1F82
		when 008067 => D <= "01110000";	-- 0x1F83
		when 008068 => D <= "01001000";	-- 0x1F84
		when 008069 => D <= "01000100";	-- 0x1F85
		when 008070 => D <= "01000010";	-- 0x1F86
		when 008071 => D <= "00000000";	-- 0x1F87
		when 008072 => D <= "00000000";	-- 0x1F88
		when 008073 => D <= "01000000";	-- 0x1F89
		when 008074 => D <= "01000000";	-- 0x1F8A
		when 008075 => D <= "01000000";	-- 0x1F8B
		when 008076 => D <= "01000000";	-- 0x1F8C
		when 008077 => D <= "01000000";	-- 0x1F8D
		when 008078 => D <= "01111110";	-- 0x1F8E
		when 008079 => D <= "00000000";	-- 0x1F8F
		when 008080 => D <= "00000000";	-- 0x1F90
		when 008081 => D <= "01000010";	-- 0x1F91
		when 008082 => D <= "01100110";	-- 0x1F92
		when 008083 => D <= "01011010";	-- 0x1F93
		when 008084 => D <= "01000010";	-- 0x1F94
		when 008085 => D <= "01000010";	-- 0x1F95
		when 008086 => D <= "01000010";	-- 0x1F96
		when 008087 => D <= "00000000";	-- 0x1F97
		when 008088 => D <= "00000000";	-- 0x1F98
		when 008089 => D <= "01000010";	-- 0x1F99
		when 008090 => D <= "01100010";	-- 0x1F9A
		when 008091 => D <= "01010010";	-- 0x1F9B
		when 008092 => D <= "01001010";	-- 0x1F9C
		when 008093 => D <= "01000110";	-- 0x1F9D
		when 008094 => D <= "01000010";	-- 0x1F9E
		when 008095 => D <= "00000000";	-- 0x1F9F
		when 008096 => D <= "00000000";	-- 0x1FA0
		when 008097 => D <= "00111100";	-- 0x1FA1
		when 008098 => D <= "01000010";	-- 0x1FA2
		when 008099 => D <= "01000010";	-- 0x1FA3
		when 008100 => D <= "01000010";	-- 0x1FA4
		when 008101 => D <= "01000010";	-- 0x1FA5
		when 008102 => D <= "00111100";	-- 0x1FA6
		when 008103 => D <= "00000000";	-- 0x1FA7
		when 008104 => D <= "00000000";	-- 0x1FA8
		when 008105 => D <= "01111100";	-- 0x1FA9
		when 008106 => D <= "01000010";	-- 0x1FAA
		when 008107 => D <= "01000010";	-- 0x1FAB
		when 008108 => D <= "01111100";	-- 0x1FAC
		when 008109 => D <= "01000000";	-- 0x1FAD
		when 008110 => D <= "01000000";	-- 0x1FAE
		when 008111 => D <= "00000000";	-- 0x1FAF
		when 008112 => D <= "00000000";	-- 0x1FB0
		when 008113 => D <= "00111100";	-- 0x1FB1
		when 008114 => D <= "01000010";	-- 0x1FB2
		when 008115 => D <= "01000010";	-- 0x1FB3
		when 008116 => D <= "01010010";	-- 0x1FB4
		when 008117 => D <= "01001010";	-- 0x1FB5
		when 008118 => D <= "00111100";	-- 0x1FB6
		when 008119 => D <= "00000000";	-- 0x1FB7
		when 008120 => D <= "00000000";	-- 0x1FB8
		when 008121 => D <= "01111100";	-- 0x1FB9
		when 008122 => D <= "01000010";	-- 0x1FBA
		when 008123 => D <= "01000010";	-- 0x1FBB
		when 008124 => D <= "01111100";	-- 0x1FBC
		when 008125 => D <= "01000100";	-- 0x1FBD
		when 008126 => D <= "01000010";	-- 0x1FBE
		when 008127 => D <= "00000000";	-- 0x1FBF
		when 008128 => D <= "00000000";	-- 0x1FC0
		when 008129 => D <= "00111100";	-- 0x1FC1
		when 008130 => D <= "01000000";	-- 0x1FC2
		when 008131 => D <= "00111100";	-- 0x1FC3
		when 008132 => D <= "00000010";	-- 0x1FC4
		when 008133 => D <= "01000010";	-- 0x1FC5
		when 008134 => D <= "00111100";	-- 0x1FC6
		when 008135 => D <= "00000000";	-- 0x1FC7
		when 008136 => D <= "00000000";	-- 0x1FC8
		when 008137 => D <= "11111110";	-- 0x1FC9
		when 008138 => D <= "00010000";	-- 0x1FCA
		when 008139 => D <= "00010000";	-- 0x1FCB
		when 008140 => D <= "00010000";	-- 0x1FCC
		when 008141 => D <= "00010000";	-- 0x1FCD
		when 008142 => D <= "00010000";	-- 0x1FCE
		when 008143 => D <= "00000000";	-- 0x1FCF
		when 008144 => D <= "00000000";	-- 0x1FD0
		when 008145 => D <= "01000010";	-- 0x1FD1
		when 008146 => D <= "01000010";	-- 0x1FD2
		when 008147 => D <= "01000010";	-- 0x1FD3
		when 008148 => D <= "01000010";	-- 0x1FD4
		when 008149 => D <= "01000010";	-- 0x1FD5
		when 008150 => D <= "00111100";	-- 0x1FD6
		when 008151 => D <= "00000000";	-- 0x1FD7
		when 008152 => D <= "00000000";	-- 0x1FD8
		when 008153 => D <= "01000010";	-- 0x1FD9
		when 008154 => D <= "01000010";	-- 0x1FDA
		when 008155 => D <= "01000010";	-- 0x1FDB
		when 008156 => D <= "01000010";	-- 0x1FDC
		when 008157 => D <= "00100100";	-- 0x1FDD
		when 008158 => D <= "00011000";	-- 0x1FDE
		when 008159 => D <= "00000000";	-- 0x1FDF
		when 008160 => D <= "00000000";	-- 0x1FE0
		when 008161 => D <= "01000010";	-- 0x1FE1
		when 008162 => D <= "01000010";	-- 0x1FE2
		when 008163 => D <= "01000010";	-- 0x1FE3
		when 008164 => D <= "01000010";	-- 0x1FE4
		when 008165 => D <= "01011010";	-- 0x1FE5
		when 008166 => D <= "00100100";	-- 0x1FE6
		when 008167 => D <= "00000000";	-- 0x1FE7
		when 008168 => D <= "00000000";	-- 0x1FE8
		when 008169 => D <= "01000010";	-- 0x1FE9
		when 008170 => D <= "00100100";	-- 0x1FEA
		when 008171 => D <= "00011000";	-- 0x1FEB
		when 008172 => D <= "00011000";	-- 0x1FEC
		when 008173 => D <= "00100100";	-- 0x1FED
		when 008174 => D <= "01000010";	-- 0x1FEE
		when 008175 => D <= "00000000";	-- 0x1FEF
		when 008176 => D <= "00000000";	-- 0x1FF0
		when 008177 => D <= "10000010";	-- 0x1FF1
		when 008178 => D <= "01000100";	-- 0x1FF2
		when 008179 => D <= "00101000";	-- 0x1FF3
		when 008180 => D <= "00010000";	-- 0x1FF4
		when 008181 => D <= "00010000";	-- 0x1FF5
		when 008182 => D <= "00010000";	-- 0x1FF6
		when 008183 => D <= "00000000";	-- 0x1FF7
		when 008184 => D <= "00000000";	-- 0x1FF8
		when 008185 => D <= "01111110";	-- 0x1FF9
		when 008186 => D <= "00000100";	-- 0x1FFA
		when 008187 => D <= "00001000";	-- 0x1FFB
		when 008188 => D <= "00010000";	-- 0x1FFC
		when 008189 => D <= "00100000";	-- 0x1FFD
		when 008190 => D <= "01111110";	-- 0x1FFE
		when 008191 => D <= "00000000";	-- 0x1FFF
		when others => D <= "--------";
		end case;
	end process;
end;
