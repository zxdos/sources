12
0e
20
4a
6f
75
73
74
20
76
32
2e
33
00
00
ff
28
f0
60
00
aa
5a
f0
55
68
00
69
03
6c
00
6d
0f
22
9e
00
e0
6a
02
7c
01
6d
07
8d
c5
4f
00
12
4e
4c
04
68
01
8b
c0
7b
01
27
48
6e
1b
6d
09
8d
c5
4f
00
12
54
fc
30
6d
3c
dd
ea
27
50
12
6a
6b
08
68
02
12
38
aa
b0
fc
33
f2
65
6d
37
f1
30
dd
ea
6d
41
f2
30
dd
ea
27
50
12
6a
6d
07
8d
c2
4d
07
19
50
28
4c
27
70
25
f8
3b
00
25
f0
6d
0f
22
9e
22
a8
46
dd
16
b0
4a
00
12
1e
22
fa
38
00
24
bc
6d
05
48
00
22
9e
6d
03
48
01
22
9e
12
80
fd
15
fd
07
3d
00
12
a0
00
ee
aa
82
f5
65
24
a0
62
00
6d
0a
ed
a1
24
9c
6d
03
ed
a1
24
90
6d
0c
ed
a1
24
96
22
ce
46
dd
00
ee
3f
00
25
16
00
ee
27
82
27
ec
8d
00
8e
10
80
24
81
34
aa
62
f5
1e
65
7f
80
52
85
40
86
00
87
10
dd
e8
aa
62
f4
1e
d0
18
41
38
66
dd
aa
82
f5
55
00
ee
4a
01
13
16
4a
02
13
0e
4a
03
13
ae
4a
04
13
b4
4a
05
13
ba
23
16
4a
02
23
68
00
ee
aa
88
f5
65
cd
03
4d
00
24
a4
23
2a
23
7a
3f
00
14
e8
00
ee
8d
60
8d
05
4f
00
8d
f7
6e
10
8e
d5
4f
00
00
ee
8d
70
8d
15
4f
00
8d
f7
6e
0c
8e
d5
4f
00
00
ee
8d
60
8d
05
4f
00
24
90
3f
00
24
96
8d
70
8d
15
3f
00
24
a0
4f
00
24
9c
91
70
24
9c
00
ee
aa
8e
f5
65
cd
01
4d
00
24
a4
23
82
3f
00
14
f0
00
ee
23
8a
aa
88
f5
55
00
ee
23
8a
aa
8e
f5
55
00
ee
27
82
27
ec
41
34
24
9c
8d
00
8e
10
80
24
81
34
aa
72
f5
1e
65
7f
80
52
85
40
dd
e8
aa
72
f4
1e
d0
18
00
ee
23
16
23
ba
00
ee
24
0e
23
ba
00
ee
aa
94
f4
65
44
02
13
ce
62
00
24
40
24
7c
aa
94
f4
55
00
ee
72
01
42
08
13
da
aa
94
f4
55
00
ee
aa
c2
d0
14
4a
04
13
ea
4a
03
14
00
6a
00
00
ee
aa
9a
f4
65
aa
94
f4
55
4b
00
6a
05
4b
00
00
ee
25
f8
6a
03
00
ee
4b
00
6a
01
4b
00
00
ee
25
f0
6a
02
00
ee
aa
9a
f4
65
44
02
14
22
62
00
24
40
24
7c
aa
9a
f4
55
00
ee
72
01
42
08
14
2e
aa
9a
f4
55
00
ee
aa
c2
d0
14
4b
00
14
3c
25
f8
6a
03
00
ee
6a
05
00
ee
41
18
14
50
41
0c
14
66
41
24
14
66
63
01
00
ee
27
ac
33
00
00
ee
6d
01
fd
18
63
fd
44
00
62
fe
44
01
62
02
00
ee
27
be
33
00
00
ee
6d
01
fd
18
63
fd
44
00
62
fe
44
01
62
02
00
ee
8d
00
8e
10
80
24
81
34
aa
c2
dd
e4
d0
14
41
38
64
02
00
ee
64
08
62
fc
00
ee
64
00
62
04
00
ee
63
fe
00
ee
63
02
00
ee
cd
01
fd
18
4d
00
24
90
4d
01
24
96
cd
01
4d
00
24
a0
4d
01
24
9c
00
ee
cd
03
3d
00
00
ee
aa
c0
f1
65
6d
3b
aa
ba
d0
d5
80
14
40
08
24
dc
40
70
24
e2
aa
c0
f1
55
00
ee
60
10
61
08
00
ee
60
68
61
f8
00
ee
24
f8
4f
00
15
92
00
ee
24
f8
4f
00
15
ce
00
ee
8d
60
8d
05
4f
00
8d
f7
6e
08
8d
e5
3f
00
00
ee
8d
70
8d
15
4f
00
8d
f7
6e
08
8d
e5
00
ee
4a
02
15
64
4a
01
15
92
4a
04
15
28
4a
05
15
3a
15
52
aa
94
f4
65
25
76
4f
00
15
46
25
84
4f
00
15
46
15
3a
27
20
27
02
27
02
aa
94
f4
65
13
da
27
20
27
02
27
02
aa
9a
f4
65
14
2e
aa
88
f5
65
25
76
4f
00
15
3a
25
84
4f
00
15
3a
15
92
aa
88
f5
65
25
76
4f
00
15
ce
25
84
4f
00
15
ce
15
92
8d
60
8d
05
4f
00
8d
f7
6e
08
8e
d5
00
ee
8d
70
8d
15
4f
00
8d
f7
6e
08
8e
d5
00
ee
aa
88
f5
65
97
10
16
62
8d
70
8d
15
3f
00
15
ec
27
0c
aa
72
f5
1e
d0
18
4a
03
15
ba
4a
02
15
c0
4a
01
6a
05
26
40
00
ee
6a
04
26
48
00
ee
26
40
aa
8e
f5
65
aa
88
f5
55
6a
03
00
ee
aa
8e
f5
65
97
10
16
78
8d
70
8d
15
3f
00
15
ec
27
0c
aa
72
f5
1e
d0
18
6a
03
26
40
00
ee
66
dd
00
ee
26
00
aa
8e
f5
55
00
ee
26
00
aa
88
f5
55
00
ee
26
1a
7b
ff
24
9c
cd
01
3d
01
24
90
3d
00
24
96
aa
72
f4
1e
d0
18
85
40
00
ee
cd
03
4d
00
16
3a
4d
01
16
34
4d
02
16
2e
60
78
61
34
00
ee
60
40
61
20
00
ee
60
40
61
08
00
ee
60
08
61
14
00
ee
26
50
aa
94
f4
55
00
ee
26
50
aa
9a
f4
55
00
ee
71
08
6d
37
8d
15
4f
00
61
37
c4
01
aa
c2
d0
14
00
ee
26
8e
3f
00
16
70
24
96
23
7a
23
7a
16
a4
24
90
23
7a
23
7a
16
98
26
8e
3f
00
16
86
24
96
23
82
23
82
16
a4
24
90
23
82
23
82
16
98
6d
03
fd
18
8d
60
8d
05
00
ee
aa
82
f5
65
24
96
22
ce
22
ce
00
ee
aa
82
f5
65
24
90
22
ce
22
ce
00
ee
27
0c
27
02
27
16
6d
0a
22
9e
79
ff
49
00
16
da
4a
01
7b
01
4a
03
7b
01
4a
02
7b
02
6a
02
4b
00
12
1e
6a
02
4b
01
6a
01
12
6a
26
e4
00
e0
27
2a
29
0c
12
12
6d
0c
fd
18
6d
18
22
9e
27
0c
27
0c
27
16
27
16
6d
20
22
9e
27
16
27
16
6d
20
22
9e
00
ee
6d
02
fd
18
6d
05
22
9e
00
ee
6d
04
fd
18
6d
0a
22
9e
00
ee
6d
08
fd
18
6d
14
22
9e
00
ee
aa
5a
f0
65
70
01
f0
55
00
ee
aa
5a
f0
65
f0
33
f2
65
6e
1b
6d
31
f0
30
dd
ea
7d
0a
f1
30
dd
ea
7d
0a
f2
30
dd
ea
00
ee
63
00
64
00
65
7c
66
3e
aa
5e
d3
43
d3
63
d5
43
d5
63
73
04
74
02
75
fc
76
fe
6d
04
22
9e
43
40
00
ee
43
80
00
ee
17
52
64
00
65
00
60
70
61
14
aa
62
d0
18
aa
82
f5
55
00
ee
41
00
17
d0
41
34
17
d8
6d
02
53
d0
17
9e
41
14
17
ac
41
08
17
be
41
20
17
be
00
ee
41
20
17
ac
41
14
17
be
41
2c
17
be
00
ee
6d
10
8d
07
4f
00
17
e8
6d
68
8d
05
4f
00
17
e8
00
ee
6d
29
8d
07
4f
00
00
ee
6d
50
8d
07
4f
00
17
e8
00
ee
6d
fe
93
d0
24
a0
00
ee
6d
02
53
d0
00
ee
48
00
17
e8
38
00
17
ac
00
ee
63
00
00
ee
42
00
00
ee
6d
04
52
d0
18
00
40
68
18
0a
40
28
18
1c
00
ee
40
10
18
0a
40
50
18
1c
00
ee
6d
11
8d
17
4f
00
00
ee
6d
21
8d
17
4f
00
18
48
00
ee
6d
1c
8d
15
4f
00
18
36
6d
05
8d
17
4f
00
00
ee
6d
15
8d
17
4f
00
18
48
00
ee
6d
1d
8d
17
4f
00
00
ee
6d
2d
8d
17
4f
00
18
48
00
ee
62
00
00
ee
00
e0
6d
00
6e
3c
aa
ac
dd
e4
6d
08
dd
e4
aa
a8
6d
10
48
00
28
a8
38
00
28
b2
aa
a8
6e
1c
6d
78
dd
e4
6d
00
dd
e4
6d
38
6e
10
dd
e4
6d
40
dd
e4
6e
28
dd
e4
6d
38
dd
e4
aa
a0
6d
48
dd
e4
6e
10
dd
e4
6d
08
6e
1c
dd
e4
aa
a4
6d
70
dd
e4
6e
28
6d
30
dd
e4
6e
10
dd
e4
28
d2
00
ee
dd
e4
7d
08
3d
80
18
a8
00
ee
6d
70
dd
e4
6d
78
dd
e4
6d
10
aa
b4
6e
3b
dd
e5
7d
08
3d
70
18
c0
60
68
61
f8
aa
c0
f1
55
00
ee
49
01
00
ee
6d
01
6e
3d
aa
5e
dd
e3
7d
04
39
02
dd
e3
7d
04
66
03
86
95
4f
00
dd
e3
00
ee
aa
c6
6d
24
6e
18
dd
e0
60
20
f0
1e
7d
10
dd
e0
f0
1e
7d
10
dd
e0
f0
1e
7d
10
dd
e0
68
00
6b
01
6a
00
25
f8
27
70
24
96
aa
82
f5
55
6d
0a
22
9e
aa
82
f5
65
29
40
22
d2
aa
82
f5
55
aa
88
f5
65
29
40
23
92
aa
88
f5
55
6d
0a
ed
9e
19
1c
00
ee
cd
0f
4d
00
24
a4
41
02
63
02
41
36
63
fe
00
ee
28
4c
27
70
aa
c2
6e
0c
6d
32
dd
e4
7d
0c
dd
e4
7d
0c
dd
e4
6e
24
6d
32
dd
e4
7d
0c
dd
e4
7d
0c
dd
e4
6e
18
6d
0a
dd
e4
6e
38
dd
e4
6d
72
dd
e4
66
00
67
00
77
01
47
6a
12
1e
6d
01
fd
18
6d
03
22
9e
aa
82
f5
65
24
a0
62
00
6d
0a
ed
a1
24
9c
6d
03
ed
a1
24
90
6d
0c
ed
a1
24
96
27
82
27
ec
8d
00
8e
10
80
24
81
34
aa
62
f5
1e
65
7f
80
52
85
40
dd
e8
aa
62
f4
1e
d0
18
41
38
1a
38
aa
82
f5
55
3f
00
29
dc
46
09
1a
48
19
84
6e
34
91
e0
19
f6
6e
14
91
e0
1a
04
6e
08
91
e0
1a
0c
6e
20
91
e0
1a
0c
00
ee
6d
70
90
d0
1a
20
6d
08
90
d0
1a
20
00
ee
6d
08
90
d0
1a
20
00
ee
6d
30
90
d0
1a
20
7d
0c
90
d0
1a
20
7d
0c
90
d0
1a
20
00
ee
7d
02
7e
04
aa
c2
dd
e4
27
02
27
02
76
01
aa
5a
f0
65
70
01
f0
55
00
ee
6d
08
fd
18
6d
14
22
9e
79
ff
49
00
16
da
12
1e
aa
5a
f0
65
70
08
f0
55
79
01
27
16
27
0c
27
16
12
1e
00
00
00
00
40
e0
40
00
66
6f
4c
ff
6c
dc
ec
78
66
f6
32
ff
36
3b
37
1e
6e
6f
4c
ff
6c
be
9e
7c
76
f6
32
ff
36
7d
79
3e
00
00
00
00
00
00
00
00
00
00
00
00
00
00
00
00
00
00
00
00
00
00
00
00
00
00
00
00
00
00
ff
ba
e8
80
ff
6d
1b
02
ff
ee
bb
b6
ff
ff
ff
ff
00
00
00
00
06
1c
28
4c
fe
00
66
24
3c
6e
00
00
00
00
60
b0
f0
60
00
c0
00
c0
00
c0
00
c0
00
c0
00
c0
00
c3
00
c7
00
cc
00
cc
c0
cc
c0
cc
c0
cc
c0
cc
7f
87
3f
03
00
00
00
00
00
00
00
00
00
00
00
00
f0
c0
f8
c0
0c
c0
0c
c0
0c
c0
0c
c0
0c
c0
0c
c0
f8
7f
f0
3f
00
00
00
00
00
00
00
00
00
00
00
00
c3
fc
c7
fc
cc
00
cc
00
c7
f0
c3
f8
c0
0c
c0
0c
cf
f8
cf
f0
00
00
00
00
30
00
30
00
30
00
30
00
fc
00
fc
00
30
00
30
00
30
00
30
00
33
00
33
00
1e
00
0c
00
