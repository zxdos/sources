6a
02
6b
0c
6c
3f
6d
0c
a2
ea
da
b6
dc
d6
6e
00
22
d4
66
03
68
02
60
60
f0
15
f0
07
30
00
12
1a
c7
17
77
08
69
ff
a2
f0
d6
71
a2
ea
da
b6
dc
d6
60
01
e0
a1
7b
fe
60
04
e0
a1
7b
02
60
1f
8b
02
da
b6
60
0c
e0
a1
7d
fe
60
0d
e0
a1
7d
02
60
1f
8d
02
dc
d6
a2
f0
d6
71
86
84
87
94
60
3f
86
02
61
1f
87
12
46
02
12
78
46
3f
12
82
47
1f
69
ff
47
00
69
01
d6
71
12
2a
68
02
63
01
80
70
80
b5
12
8a
68
fe
63
0a
80
70
80
d5
3f
01
12
a2
61
02
80
15
3f
01
12
ba
80
15
3f
01
12
c8
80
15
3f
01
12
c2
60
20
f0
18
22
d4
8e
34
22
d4
66
3e
33
01
66
03
68
fe
33
01
68
02
12
16
79
ff
49
fe
69
ff
12
c8
79
01
49
02
69
01
60
04
f0
18
76
01
46
40
76
fe
12
6c
a2
f2
fe
33
f2
65
f1
29
64
14
65
00
d4
55
74
15
f2
29
d4
55
00
ee
80
80
80
80
80
80
80
00
00
00
00
00
