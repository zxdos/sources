-- ZPU
--
-- Copyright 2004-2008 oharboe - �yvind Harboe - oyvind.harboe@zylin.com
-- Modified by Alastair M. Robinson for the ZPUFlex project.
--
-- The FreeBSD license
-- 
-- Redistribution and use in source and binary forms, with or without
-- modification, are permitted provided that the following conditions
-- are met:
-- 
-- 1. Redistributions of source code must retain the above copyright
--    notice, this list of conditions and the following disclaimer.
-- 2. Redistributions in binary form must reproduce the above
--    copyright notice, this list of conditions and the following
--    disclaimer in the documentation and/or other materials
--    provided with the distribution.
-- 
-- THIS SOFTWARE IS PROVIDED BY THE ZPU PROJECT ``AS IS'' AND ANY
-- EXPRESS OR IMPLIED WARRANTIES, INCLUDING, BUT NOT LIMITED TO,
-- THE IMPLIED WARRANTIES OF MERCHANTABILITY AND FITNESS FOR A
-- PARTICULAR PURPOSE ARE DISCLAIMED. IN NO EVENT SHALL THE
-- ZPU PROJECT OR CONTRIBUTORS BE LIABLE FOR ANY DIRECT,
-- INDIRECT, INCIDENTAL, SPECIAL, EXEMPLARY, OR CONSEQUENTIAL DAMAGES
-- (INCLUDING, BUT NOT LIMITED TO, PROCUREMENT OF SUBSTITUTE GOODS
-- OR SERVICES; LOSS OF USE, DATA, OR PROFITS; OR BUSINESS INTERRUPTION)
-- HOWEVER CAUSED AND ON ANY THEORY OF LIABILITY, WHETHER IN CONTRACT,
-- STRICT LIABILITY, OR TORT (INCLUDING NEGLIGENCE OR OTHERWISE)
-- ARISING IN ANY WAY OUT OF THE USE OF THIS SOFTWARE, EVEN IF
-- ADVISED OF THE POSSIBILITY OF SUCH DAMAGE.
-- 
-- The views and conclusions contained in the software and documentation
-- are those of the authors and should not be interpreted as representing
-- official policies, either expressed or implied, of the ZPU Project.

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;


library work;
use work.zpupkg.all;

entity CtrlROM_ROM is
generic
	(
		maxAddrBitBRAM : integer := maxAddrBitBRAMLimit -- Specify your actual ROM size to save LEs and unnecessary block RAM usage.
	);
port (
	clk : in std_logic;
	areset : in std_logic := '0';
	from_zpu : in ZPU_ToROM;
	to_zpu : out ZPU_FromROM
);
end CtrlROM_ROM;

architecture arch of CtrlROM_ROM is

type ram_type is array(natural range 0 to ((2**(maxAddrBitBRAM+1))/4)-1) of std_logic_vector(wordSize-1 downto 0);

shared variable ram : ram_type :=
(
     0 => x"0b0b0b0b",
     1 => x"8c0b0b0b",
     2 => x"0b81e004",
     3 => x"0b0b0b0b",
     4 => x"8c04ff0d",
     5 => x"80040400",
     6 => x"00000016",
     7 => x"00000000",
     8 => x"0b0b80c8",
     9 => x"b4080b0b",
    10 => x"80c8b808",
    11 => x"0b0b80c8",
    12 => x"bc080b0b",
    13 => x"0b0b9808",
    14 => x"2d0b0b80",
    15 => x"c8bc0c0b",
    16 => x"0b80c8b8",
    17 => x"0c0b0b80",
    18 => x"c8b40c04",
    19 => x"00000000",
    20 => x"00000000",
    21 => x"00000000",
    22 => x"00000000",
    23 => x"00000000",
    24 => x"71fd0608",
    25 => x"72830609",
    26 => x"81058205",
    27 => x"832b2a83",
    28 => x"ffff0652",
    29 => x"0471fc06",
    30 => x"08728306",
    31 => x"09810583",
    32 => x"05101010",
    33 => x"2a81ff06",
    34 => x"520471fd",
    35 => x"060883ff",
    36 => x"ff738306",
    37 => x"09810582",
    38 => x"05832b2b",
    39 => x"09067383",
    40 => x"ffff0673",
    41 => x"83060981",
    42 => x"05820583",
    43 => x"2b0b2b07",
    44 => x"72fc060c",
    45 => x"51510471",
    46 => x"fc06080b",
    47 => x"0b0bbab8",
    48 => x"73830610",
    49 => x"10050806",
    50 => x"7381ff06",
    51 => x"73830609",
    52 => x"81058305",
    53 => x"1010102b",
    54 => x"0772fc06",
    55 => x"0c515104",
    56 => x"80c8b470",
    57 => x"80d2f427",
    58 => x"8b388071",
    59 => x"70840553",
    60 => x"0c81e304",
    61 => x"8c518a83",
    62 => x"0402fc05",
    63 => x"0df88051",
    64 => x"8f0b80c8",
    65 => x"c40c9f0b",
    66 => x"80c8c80c",
    67 => x"a0717081",
    68 => x"05533480",
    69 => x"c8c808ff",
    70 => x"0580c8c8",
    71 => x"0c80c8c8",
    72 => x"088025e8",
    73 => x"3880c8c4",
    74 => x"08ff0580",
    75 => x"c8c40c80",
    76 => x"c8c40880",
    77 => x"25d03880",
    78 => x"0b80c8c8",
    79 => x"0c800b80",
    80 => x"c8c40c02",
    81 => x"84050d04",
    82 => x"02f0050d",
    83 => x"f88053f8",
    84 => x"a05483bf",
    85 => x"52737081",
    86 => x"05553351",
    87 => x"70737081",
    88 => x"055534ff",
    89 => x"12527180",
    90 => x"25eb38fb",
    91 => x"c0539f52",
    92 => x"a0737081",
    93 => x"055534ff",
    94 => x"12527180",
    95 => x"25f23802",
    96 => x"90050d04",
    97 => x"02f4050d",
    98 => x"74538e0b",
    99 => x"80c8c408",
   100 => x"25913882",
   101 => x"c82d80c8",
   102 => x"c408ff05",
   103 => x"80c8c40c",
   104 => x"838a0480",
   105 => x"c8c40880",
   106 => x"c8c80853",
   107 => x"51728a2e",
   108 => x"098106be",
   109 => x"38715171",
   110 => x"9f24a438",
   111 => x"80c8c408",
   112 => x"a02911f8",
   113 => x"80115151",
   114 => x"a0713480",
   115 => x"c8c80881",
   116 => x"0580c8c8",
   117 => x"0c80c8c8",
   118 => x"08519f71",
   119 => x"25de3880",
   120 => x"0b80c8c8",
   121 => x"0c80c8c4",
   122 => x"08810580",
   123 => x"c8c40c84",
   124 => x"880470a0",
   125 => x"2912f880",
   126 => x"11515172",
   127 => x"713480c8",
   128 => x"c8088105",
   129 => x"80c8c80c",
   130 => x"80c8c808",
   131 => x"a02e0981",
   132 => x"06913880",
   133 => x"0b80c8c8",
   134 => x"0c80c8c4",
   135 => x"08810580",
   136 => x"c8c40c02",
   137 => x"8c050d04",
   138 => x"02e8050d",
   139 => x"77795656",
   140 => x"880bfc16",
   141 => x"77712c8f",
   142 => x"06545254",
   143 => x"80537272",
   144 => x"25953871",
   145 => x"53fbe014",
   146 => x"51877134",
   147 => x"8114ff14",
   148 => x"545472f1",
   149 => x"387153f9",
   150 => x"1576712c",
   151 => x"87065351",
   152 => x"71802e8b",
   153 => x"38fbe014",
   154 => x"51717134",
   155 => x"81145472",
   156 => x"8e249538",
   157 => x"8f733153",
   158 => x"fbe01451",
   159 => x"a0713481",
   160 => x"14ff1454",
   161 => x"5472f138",
   162 => x"0298050d",
   163 => x"0402ec05",
   164 => x"0d800b80",
   165 => x"c8cc0cf6",
   166 => x"8c08f690",
   167 => x"0871882c",
   168 => x"565381ff",
   169 => x"06537373",
   170 => x"25893872",
   171 => x"54820b80",
   172 => x"c8cc0c71",
   173 => x"882c7281",
   174 => x"ff065355",
   175 => x"7472258d",
   176 => x"387180c8",
   177 => x"cc088407",
   178 => x"80c8cc0c",
   179 => x"5573842b",
   180 => x"75832b56",
   181 => x"5485bc74",
   182 => x"258f3882",
   183 => x"0b0b0b80",
   184 => x"c19c0c80",
   185 => x"d05385f3",
   186 => x"04810b0b",
   187 => x"0b80c19c",
   188 => x"0cbc530b",
   189 => x"0b80c19c",
   190 => x"0881712b",
   191 => x"ff05f688",
   192 => x"0cfc0875",
   193 => x"7531ffb0",
   194 => x"05ff1371",
   195 => x"712cff94",
   196 => x"1a709f2a",
   197 => x"1170812c",
   198 => x"80c8cc08",
   199 => x"52545153",
   200 => x"57535152",
   201 => x"5276802e",
   202 => x"85387081",
   203 => x"075170f6",
   204 => x"940c7209",
   205 => x"8105f680",
   206 => x"0c710981",
   207 => x"05f6840c",
   208 => x"0294050d",
   209 => x"0402f405",
   210 => x"0d745372",
   211 => x"70810554",
   212 => x"80f52d52",
   213 => x"71802e89",
   214 => x"38715183",
   215 => x"842d86cb",
   216 => x"04810b80",
   217 => x"c8b40c02",
   218 => x"8c050d04",
   219 => x"02fc050d",
   220 => x"81808051",
   221 => x"c0115170",
   222 => x"fb380284",
   223 => x"050d0402",
   224 => x"fc050dec",
   225 => x"5183710c",
   226 => x"86ec2d82",
   227 => x"710c0284",
   228 => x"050d0402",
   229 => x"fc050d84",
   230 => x"bf5186ec",
   231 => x"2dff1151",
   232 => x"708025f6",
   233 => x"38028405",
   234 => x"0d040402",
   235 => x"fc050d8f",
   236 => x"f12d80c8",
   237 => x"b40880c5",
   238 => x"f00c80c4",
   239 => x"d85192a6",
   240 => x"2d028405",
   241 => x"0d0402fc",
   242 => x"050d8ff1",
   243 => x"2d80c8b4",
   244 => x"0880c4c8",
   245 => x"0c80c3b0",
   246 => x"5192a62d",
   247 => x"0284050d",
   248 => x"0402dc05",
   249 => x"0d7a5480",
   250 => x"59840bec",
   251 => x"0c80c8dc",
   252 => x"08828007",
   253 => x"82803270",
   254 => x"80c8dc0c",
   255 => x"fc0c86ec",
   256 => x"2d735280",
   257 => x"c8d051b1",
   258 => x"9c2d80c8",
   259 => x"b408792e",
   260 => x"81ac3880",
   261 => x"c8d40855",
   262 => x"74852e09",
   263 => x"8106a538",
   264 => x"735186c5",
   265 => x"2d87932d",
   266 => x"87932d87",
   267 => x"932d8793",
   268 => x"2d87932d",
   269 => x"87932d80",
   270 => x"c8e00851",
   271 => x"92a62d81",
   272 => x"5389f904",
   273 => x"74f80ca5",
   274 => x"0bec0c87",
   275 => x"932d840b",
   276 => x"ec0c78ff",
   277 => x"16555873",
   278 => x"802e8b38",
   279 => x"81187481",
   280 => x"2a555888",
   281 => x"d704f718",
   282 => x"58815980",
   283 => x"752580ce",
   284 => x"38775273",
   285 => x"5184a82d",
   286 => x"80c9ac52",
   287 => x"80c8d051",
   288 => x"b3e92d80",
   289 => x"c8b40880",
   290 => x"2e9b3880",
   291 => x"c9ac5783",
   292 => x"fc567670",
   293 => x"84055808",
   294 => x"e80cfc16",
   295 => x"56758025",
   296 => x"f13889ad",
   297 => x"0480c8b4",
   298 => x"08598480",
   299 => x"5580c8d0",
   300 => x"51b3b92d",
   301 => x"fc801581",
   302 => x"15555588",
   303 => x"eb04800b",
   304 => x"80c1a00c",
   305 => x"80c8dc08",
   306 => x"82800782",
   307 => x"80327080",
   308 => x"c8dc0cfc",
   309 => x"0c78802e",
   310 => x"973880c8",
   311 => x"e0085192",
   312 => x"a62d810b",
   313 => x"ec0c8793",
   314 => x"2d820bec",
   315 => x"0c89f704",
   316 => x"80c38c51",
   317 => x"92a62d78",
   318 => x"537280c8",
   319 => x"b40c02a4",
   320 => x"050d0402",
   321 => x"f4050d84",
   322 => x"0b80c8dc",
   323 => x"0c805186",
   324 => x"ff2d840b",
   325 => x"ec0c8fc1",
   326 => x"2d8bec2d",
   327 => x"81f92d83",
   328 => x"528fa42d",
   329 => x"8151858d",
   330 => x"2dff1252",
   331 => x"718025f1",
   332 => x"38840bec",
   333 => x"0cbfd051",
   334 => x"86c52da7",
   335 => x"d42d80c8",
   336 => x"b408802e",
   337 => x"818f3881",
   338 => x"0bec0c84",
   339 => x"0bec0c87",
   340 => x"e151bab1",
   341 => x"2d80c8dc",
   342 => x"0870822c",
   343 => x"80c6c80c",
   344 => x"fc0c80c9",
   345 => x"8c08882a",
   346 => x"70810651",
   347 => x"5271802e",
   348 => x"8c3880c2",
   349 => x"a00b80c8",
   350 => x"e00c8b85",
   351 => x"0480c1a4",
   352 => x"0b80c8e0",
   353 => x"0c80c8e0",
   354 => x"085192a6",
   355 => x"2d840b80",
   356 => x"c9a00c8f",
   357 => x"fa2d8bf8",
   358 => x"2d92b92d",
   359 => x"80c8e008",
   360 => x"ac1180f5",
   361 => x"2d7080c8",
   362 => x"dc0c80c6",
   363 => x"c8088106",
   364 => x"52545271",
   365 => x"802e8838",
   366 => x"72840780",
   367 => x"c8dc0c80",
   368 => x"c8dc08fc",
   369 => x"0c865280",
   370 => x"c8b40883",
   371 => x"38845271",
   372 => x"ec0c8b96",
   373 => x"04800b80",
   374 => x"c8b40c02",
   375 => x"8c050d04",
   376 => x"71980c04",
   377 => x"ffb00880",
   378 => x"c8b40c04",
   379 => x"810bffb0",
   380 => x"0c04800b",
   381 => x"ffb00c04",
   382 => x"02f4050d",
   383 => x"8d860480",
   384 => x"c8b40881",
   385 => x"f02e0981",
   386 => x"068a3881",
   387 => x"0b80c6c0",
   388 => x"0c8d8604",
   389 => x"80c8b408",
   390 => x"81e02e09",
   391 => x"81068a38",
   392 => x"810b80c6",
   393 => x"c40c8d86",
   394 => x"0480c8b4",
   395 => x"085280c6",
   396 => x"c408802e",
   397 => x"893880c8",
   398 => x"b4088180",
   399 => x"05527184",
   400 => x"2c728f06",
   401 => x"535380c6",
   402 => x"c008802e",
   403 => x"9a387284",
   404 => x"2980c680",
   405 => x"05721381",
   406 => x"712b7009",
   407 => x"73080673",
   408 => x"0c515353",
   409 => x"8cfa0472",
   410 => x"842980c6",
   411 => x"80057213",
   412 => x"83712b72",
   413 => x"0807720c",
   414 => x"5353800b",
   415 => x"80c6c40c",
   416 => x"800b80c6",
   417 => x"c00c80c8",
   418 => x"e4518e8d",
   419 => x"2d80c8b4",
   420 => x"08ff24fe",
   421 => x"ea38800b",
   422 => x"80c8b40c",
   423 => x"028c050d",
   424 => x"0402f805",
   425 => x"0d80c680",
   426 => x"528f5180",
   427 => x"72708405",
   428 => x"540cff11",
   429 => x"51708025",
   430 => x"f2380288",
   431 => x"050d0402",
   432 => x"f0050d75",
   433 => x"518bf22d",
   434 => x"70822cfc",
   435 => x"0680c680",
   436 => x"1172109e",
   437 => x"06710870",
   438 => x"722a7083",
   439 => x"0682742b",
   440 => x"70097406",
   441 => x"760c5451",
   442 => x"56575351",
   443 => x"538bec2d",
   444 => x"7180c8b4",
   445 => x"0c029005",
   446 => x"0d0402fc",
   447 => x"050d7251",
   448 => x"80710c80",
   449 => x"0b84120c",
   450 => x"0284050d",
   451 => x"0402f005",
   452 => x"0d757008",
   453 => x"84120853",
   454 => x"5353ff54",
   455 => x"71712ea8",
   456 => x"388bf22d",
   457 => x"84130870",
   458 => x"84291488",
   459 => x"11700870",
   460 => x"81ff0684",
   461 => x"18088111",
   462 => x"8706841a",
   463 => x"0c535155",
   464 => x"5151518b",
   465 => x"ec2d7154",
   466 => x"7380c8b4",
   467 => x"0c029005",
   468 => x"0d0402f4",
   469 => x"050d8bf2",
   470 => x"2de00870",
   471 => x"8b2a7081",
   472 => x"06515253",
   473 => x"70802ea1",
   474 => x"3880c8e4",
   475 => x"08708429",
   476 => x"80c8ec05",
   477 => x"7481ff06",
   478 => x"710c5151",
   479 => x"80c8e408",
   480 => x"81118706",
   481 => x"80c8e40c",
   482 => x"51728c2c",
   483 => x"83ff0680",
   484 => x"c98c0c80",
   485 => x"0b80c990",
   486 => x"0c8be42d",
   487 => x"8bec2d02",
   488 => x"8c050d04",
   489 => x"02fc050d",
   490 => x"8bf22d81",
   491 => x"0b80c990",
   492 => x"0c8bec2d",
   493 => x"80c99008",
   494 => x"5170f938",
   495 => x"0284050d",
   496 => x"0402fc05",
   497 => x"0d80c8e4",
   498 => x"518dfa2d",
   499 => x"8da12d8e",
   500 => x"d2518be0",
   501 => x"2d028405",
   502 => x"0d0402fc",
   503 => x"050d8fcf",
   504 => x"5186ec2d",
   505 => x"ff115170",
   506 => x"8025f638",
   507 => x"0284050d",
   508 => x"0480c998",
   509 => x"0880c8b4",
   510 => x"0c0402fc",
   511 => x"050d810b",
   512 => x"80c6f40c",
   513 => x"8151858d",
   514 => x"2d028405",
   515 => x"0d0402fc",
   516 => x"050d9098",
   517 => x"048bf82d",
   518 => x"80f6518d",
   519 => x"bf2d80c8",
   520 => x"b408f238",
   521 => x"80da518d",
   522 => x"bf2d80c8",
   523 => x"b408e638",
   524 => x"80c6f008",
   525 => x"518dbf2d",
   526 => x"80c8b408",
   527 => x"d83880c8",
   528 => x"b40880c6",
   529 => x"f40c80c8",
   530 => x"b4085185",
   531 => x"8d2d0284",
   532 => x"050d0402",
   533 => x"ec050d76",
   534 => x"54805287",
   535 => x"0b881580",
   536 => x"f52d5653",
   537 => x"74722483",
   538 => x"38a05372",
   539 => x"5183842d",
   540 => x"81128b15",
   541 => x"80f52d54",
   542 => x"52727225",
   543 => x"de380294",
   544 => x"050d0402",
   545 => x"f0050d80",
   546 => x"c9980854",
   547 => x"81f92d80",
   548 => x"0b80c99c",
   549 => x"0c730880",
   550 => x"2e818638",
   551 => x"820b80c8",
   552 => x"c80c80c9",
   553 => x"9c088f06",
   554 => x"80c8c40c",
   555 => x"73085271",
   556 => x"832e9638",
   557 => x"71832689",
   558 => x"3871812e",
   559 => x"af38928a",
   560 => x"0471852e",
   561 => x"9f38928a",
   562 => x"04881480",
   563 => x"f52d8415",
   564 => x"08bfe853",
   565 => x"545286c5",
   566 => x"2d718429",
   567 => x"13700852",
   568 => x"52928e04",
   569 => x"735190d3",
   570 => x"2d928a04",
   571 => x"80c6c808",
   572 => x"8815082c",
   573 => x"70810651",
   574 => x"5271802e",
   575 => x"8738bfec",
   576 => x"51928704",
   577 => x"bff05186",
   578 => x"c52d8414",
   579 => x"085186c5",
   580 => x"2d80c99c",
   581 => x"08810580",
   582 => x"c99c0c8c",
   583 => x"14549195",
   584 => x"04029005",
   585 => x"0d047180",
   586 => x"c9980c91",
   587 => x"832d80c9",
   588 => x"9c08ff05",
   589 => x"80c9a00c",
   590 => x"0402e805",
   591 => x"0d80c998",
   592 => x"0880c9a4",
   593 => x"08575580",
   594 => x"f6518dbf",
   595 => x"2d80c8b4",
   596 => x"08812a70",
   597 => x"81065152",
   598 => x"71802ea2",
   599 => x"3892e304",
   600 => x"8bf82d80",
   601 => x"f6518dbf",
   602 => x"2d80c8b4",
   603 => x"08f23880",
   604 => x"c6f40881",
   605 => x"327080c6",
   606 => x"f40c5185",
   607 => x"8d2d800b",
   608 => x"80c9940c",
   609 => x"86518dbf",
   610 => x"2d80c8b4",
   611 => x"08812a70",
   612 => x"81065152",
   613 => x"71802e8b",
   614 => x"3880c8dc",
   615 => x"08903280",
   616 => x"c8dc0c8c",
   617 => x"518dbf2d",
   618 => x"80c8b408",
   619 => x"812a7081",
   620 => x"06515271",
   621 => x"802e80d1",
   622 => x"3880c6cc",
   623 => x"0880c6e0",
   624 => x"0880c6cc",
   625 => x"0c80c6e0",
   626 => x"0c80c6d0",
   627 => x"0880c6e4",
   628 => x"0880c6d0",
   629 => x"0c80c6e4",
   630 => x"0c80c6d4",
   631 => x"0880c6e8",
   632 => x"0880c6d4",
   633 => x"0c80c6e8",
   634 => x"0c80c6d8",
   635 => x"0880c6ec",
   636 => x"0880c6d8",
   637 => x"0c80c6ec",
   638 => x"0c80c6dc",
   639 => x"0880c6f0",
   640 => x"0880c6dc",
   641 => x"0c80c6f0",
   642 => x"0c80c98c",
   643 => x"08a00652",
   644 => x"80722596",
   645 => x"388fda2d",
   646 => x"8bf82d80",
   647 => x"c6f40881",
   648 => x"327080c6",
   649 => x"f40c5185",
   650 => x"8d2d80c6",
   651 => x"f40882ef",
   652 => x"3880c6e0",
   653 => x"08518dbf",
   654 => x"2d80c8b4",
   655 => x"08802e8b",
   656 => x"3880c994",
   657 => x"08810780",
   658 => x"c9940c80",
   659 => x"c6e40851",
   660 => x"8dbf2d80",
   661 => x"c8b40880",
   662 => x"2e8b3880",
   663 => x"c9940882",
   664 => x"0780c994",
   665 => x"0c80c6e8",
   666 => x"08518dbf",
   667 => x"2d80c8b4",
   668 => x"08802e8b",
   669 => x"3880c994",
   670 => x"08840780",
   671 => x"c9940c80",
   672 => x"c6ec0851",
   673 => x"8dbf2d80",
   674 => x"c8b40880",
   675 => x"2e8b3880",
   676 => x"c9940888",
   677 => x"0780c994",
   678 => x"0c80c6f0",
   679 => x"08518dbf",
   680 => x"2d80c8b4",
   681 => x"08802e8b",
   682 => x"3880c994",
   683 => x"08900780",
   684 => x"c9940c80",
   685 => x"c6cc0851",
   686 => x"8dbf2d80",
   687 => x"c8b40880",
   688 => x"2e8c3880",
   689 => x"c9940882",
   690 => x"800780c9",
   691 => x"940c80c6",
   692 => x"d008518d",
   693 => x"bf2d80c8",
   694 => x"b408802e",
   695 => x"8c3880c9",
   696 => x"94088480",
   697 => x"0780c994",
   698 => x"0c80c6d4",
   699 => x"08518dbf",
   700 => x"2d80c8b4",
   701 => x"08802e8c",
   702 => x"3880c994",
   703 => x"08888007",
   704 => x"80c9940c",
   705 => x"80c6d808",
   706 => x"518dbf2d",
   707 => x"80c8b408",
   708 => x"802e8c38",
   709 => x"80c99408",
   710 => x"90800780",
   711 => x"c9940c80",
   712 => x"c6dc0851",
   713 => x"8dbf2d80",
   714 => x"c8b40880",
   715 => x"2e8c3880",
   716 => x"c99408a0",
   717 => x"800780c9",
   718 => x"940c9451",
   719 => x"8dbf2d80",
   720 => x"c8b40852",
   721 => x"91518dbf",
   722 => x"2d7180c8",
   723 => x"b4080652",
   724 => x"80e6518d",
   725 => x"bf2d7180",
   726 => x"c8b40806",
   727 => x"5271802e",
   728 => x"8d3880c9",
   729 => x"94088480",
   730 => x"800780c9",
   731 => x"940c80fe",
   732 => x"518dbf2d",
   733 => x"80c8b408",
   734 => x"5287518d",
   735 => x"bf2d7180",
   736 => x"c8b40807",
   737 => x"5271802e",
   738 => x"8d3880c9",
   739 => x"94088880",
   740 => x"800780c9",
   741 => x"940c80c9",
   742 => x"9408ed0c",
   743 => x"9faa0494",
   744 => x"518dbf2d",
   745 => x"80c8b408",
   746 => x"5291518d",
   747 => x"bf2d7180",
   748 => x"c8b40806",
   749 => x"5280e651",
   750 => x"8dbf2d71",
   751 => x"80c8b408",
   752 => x"06527180",
   753 => x"2e8d3880",
   754 => x"c9940884",
   755 => x"80800780",
   756 => x"c9940c80",
   757 => x"fe518dbf",
   758 => x"2d80c8b4",
   759 => x"08528751",
   760 => x"8dbf2d71",
   761 => x"80c8b408",
   762 => x"07527180",
   763 => x"2e8d3880",
   764 => x"c9940888",
   765 => x"80800780",
   766 => x"c9940c80",
   767 => x"c99408ed",
   768 => x"0c81f551",
   769 => x"8dbf2d80",
   770 => x"c8b40881",
   771 => x"2a708106",
   772 => x"515271a4",
   773 => x"3880c6e0",
   774 => x"08518dbf",
   775 => x"2d80c8b4",
   776 => x"08812a70",
   777 => x"81065152",
   778 => x"718e3880",
   779 => x"c98c0881",
   780 => x"06528072",
   781 => x"2580c238",
   782 => x"80c98c08",
   783 => x"81065280",
   784 => x"72258438",
   785 => x"8fda2d80",
   786 => x"c9a00852",
   787 => x"71802e8a",
   788 => x"38ff1280",
   789 => x"c9a00c98",
   790 => x"f90480c9",
   791 => x"9c081080",
   792 => x"c99c0805",
   793 => x"70842916",
   794 => x"51528812",
   795 => x"08802e89",
   796 => x"38ff5188",
   797 => x"12085271",
   798 => x"2d81f251",
   799 => x"8dbf2d80",
   800 => x"c8b40881",
   801 => x"2a708106",
   802 => x"515271a4",
   803 => x"3880c6e4",
   804 => x"08518dbf",
   805 => x"2d80c8b4",
   806 => x"08812a70",
   807 => x"81065152",
   808 => x"718e3880",
   809 => x"c98c0882",
   810 => x"06528072",
   811 => x"2580c338",
   812 => x"80c98c08",
   813 => x"82065280",
   814 => x"72258438",
   815 => x"8fda2d80",
   816 => x"c99c08ff",
   817 => x"1180c9a0",
   818 => x"08565353",
   819 => x"7372258a",
   820 => x"38811480",
   821 => x"c9a00c99",
   822 => x"f2047210",
   823 => x"13708429",
   824 => x"16515288",
   825 => x"1208802e",
   826 => x"8938fe51",
   827 => x"88120852",
   828 => x"712d81fd",
   829 => x"518dbf2d",
   830 => x"80c8b408",
   831 => x"812a7081",
   832 => x"06515271",
   833 => x"a43880c6",
   834 => x"e808518d",
   835 => x"bf2d80c8",
   836 => x"b408812a",
   837 => x"70810651",
   838 => x"52718e38",
   839 => x"80c98c08",
   840 => x"84065280",
   841 => x"722580c0",
   842 => x"3880c98c",
   843 => x"08840652",
   844 => x"80722584",
   845 => x"388fda2d",
   846 => x"80c9a008",
   847 => x"802e8a38",
   848 => x"800b80c9",
   849 => x"a00c9ae8",
   850 => x"0480c99c",
   851 => x"081080c9",
   852 => x"9c080570",
   853 => x"84291651",
   854 => x"52881208",
   855 => x"802e8938",
   856 => x"fd518812",
   857 => x"0852712d",
   858 => x"81fa518d",
   859 => x"bf2d80c8",
   860 => x"b408812a",
   861 => x"70810651",
   862 => x"5271a438",
   863 => x"80c6ec08",
   864 => x"518dbf2d",
   865 => x"80c8b408",
   866 => x"812a7081",
   867 => x"06515271",
   868 => x"8e3880c9",
   869 => x"8c088806",
   870 => x"52807225",
   871 => x"80c03880",
   872 => x"c98c0888",
   873 => x"06528072",
   874 => x"2584388f",
   875 => x"da2d80c9",
   876 => x"9c08ff11",
   877 => x"545280c9",
   878 => x"a0087325",
   879 => x"89387280",
   880 => x"c9a00c9b",
   881 => x"de047110",
   882 => x"12708429",
   883 => x"16515288",
   884 => x"1208802e",
   885 => x"8938fc51",
   886 => x"88120852",
   887 => x"712d80c9",
   888 => x"a0087053",
   889 => x"5473802e",
   890 => x"8a388c15",
   891 => x"ff155555",
   892 => x"9be50482",
   893 => x"0b80c8c8",
   894 => x"0c718f06",
   895 => x"80c8c40c",
   896 => x"81eb518d",
   897 => x"bf2d80c8",
   898 => x"b408812a",
   899 => x"70810651",
   900 => x"5271802e",
   901 => x"ad387408",
   902 => x"852e0981",
   903 => x"06a43888",
   904 => x"1580f52d",
   905 => x"ff055271",
   906 => x"881681b7",
   907 => x"2d71982b",
   908 => x"52718025",
   909 => x"8838800b",
   910 => x"881681b7",
   911 => x"2d745190",
   912 => x"d32d81f4",
   913 => x"518dbf2d",
   914 => x"80c8b408",
   915 => x"812a7081",
   916 => x"06515271",
   917 => x"802eb338",
   918 => x"7408852e",
   919 => x"098106aa",
   920 => x"38881580",
   921 => x"f52d8105",
   922 => x"52718816",
   923 => x"81b72d71",
   924 => x"81ff068b",
   925 => x"1680f52d",
   926 => x"54527272",
   927 => x"27873872",
   928 => x"881681b7",
   929 => x"2d745190",
   930 => x"d32d80da",
   931 => x"518dbf2d",
   932 => x"80c8b408",
   933 => x"812a7081",
   934 => x"06515271",
   935 => x"8e3880c9",
   936 => x"8c089006",
   937 => x"52807225",
   938 => x"81bc3880",
   939 => x"c9980880",
   940 => x"c98c0890",
   941 => x"06535380",
   942 => x"72258438",
   943 => x"8fda2d80",
   944 => x"c9a00854",
   945 => x"73802e8a",
   946 => x"388c13ff",
   947 => x"1555539d",
   948 => x"c4047208",
   949 => x"5271822e",
   950 => x"a6387182",
   951 => x"26893871",
   952 => x"812eaa38",
   953 => x"9ee60471",
   954 => x"832eb438",
   955 => x"71842e09",
   956 => x"810680f2",
   957 => x"38881308",
   958 => x"5192a62d",
   959 => x"9ee60480",
   960 => x"c9a00851",
   961 => x"88130852",
   962 => x"712d9ee6",
   963 => x"04810b88",
   964 => x"14082b80",
   965 => x"c6c80832",
   966 => x"80c6c80c",
   967 => x"9eba0488",
   968 => x"1380f52d",
   969 => x"81058b14",
   970 => x"80f52d53",
   971 => x"54717424",
   972 => x"83388054",
   973 => x"73881481",
   974 => x"b72d9183",
   975 => x"2d9ee604",
   976 => x"7508802e",
   977 => x"a4387508",
   978 => x"518dbf2d",
   979 => x"80c8b408",
   980 => x"81065271",
   981 => x"802e8c38",
   982 => x"80c9a008",
   983 => x"51841608",
   984 => x"52712d88",
   985 => x"165675d8",
   986 => x"38805480",
   987 => x"0b80c8c8",
   988 => x"0c738f06",
   989 => x"80c8c40c",
   990 => x"a0527380",
   991 => x"c9a0082e",
   992 => x"09810699",
   993 => x"3880c99c",
   994 => x"08ff0574",
   995 => x"32700981",
   996 => x"05707207",
   997 => x"9f2a9171",
   998 => x"31515153",
   999 => x"53715183",
  1000 => x"842d8114",
  1001 => x"548e7425",
  1002 => x"c23880c6",
  1003 => x"f40880c8",
  1004 => x"b40c0298",
  1005 => x"050d0402",
  1006 => x"f4050dd4",
  1007 => x"5281ff72",
  1008 => x"0c710853",
  1009 => x"81ff720c",
  1010 => x"72882b83",
  1011 => x"fe800672",
  1012 => x"087081ff",
  1013 => x"06515253",
  1014 => x"81ff720c",
  1015 => x"72710788",
  1016 => x"2b720870",
  1017 => x"81ff0651",
  1018 => x"525381ff",
  1019 => x"720c7271",
  1020 => x"07882b72",
  1021 => x"087081ff",
  1022 => x"06720780",
  1023 => x"c8b40c52",
  1024 => x"53028c05",
  1025 => x"0d0402f4",
  1026 => x"050d7476",
  1027 => x"7181ff06",
  1028 => x"d40c5353",
  1029 => x"80c9a808",
  1030 => x"85387189",
  1031 => x"2b527198",
  1032 => x"2ad40c71",
  1033 => x"902a7081",
  1034 => x"ff06d40c",
  1035 => x"5171882a",
  1036 => x"7081ff06",
  1037 => x"d40c5171",
  1038 => x"81ff06d4",
  1039 => x"0c72902a",
  1040 => x"7081ff06",
  1041 => x"d40c51d4",
  1042 => x"087081ff",
  1043 => x"06515182",
  1044 => x"b8bf5270",
  1045 => x"81ff2e09",
  1046 => x"81069438",
  1047 => x"81ff0bd4",
  1048 => x"0cd40870",
  1049 => x"81ff06ff",
  1050 => x"14545151",
  1051 => x"71e53870",
  1052 => x"80c8b40c",
  1053 => x"028c050d",
  1054 => x"0402fc05",
  1055 => x"0d81c751",
  1056 => x"81ff0bd4",
  1057 => x"0cff1151",
  1058 => x"708025f4",
  1059 => x"38028405",
  1060 => x"0d0402f4",
  1061 => x"050d81ff",
  1062 => x"0bd40c93",
  1063 => x"53805287",
  1064 => x"fc80c151",
  1065 => x"a0862d80",
  1066 => x"c8b4088b",
  1067 => x"3881ff0b",
  1068 => x"d40c8153",
  1069 => x"a1c004a0",
  1070 => x"f92dff13",
  1071 => x"5372de38",
  1072 => x"7280c8b4",
  1073 => x"0c028c05",
  1074 => x"0d0402ec",
  1075 => x"050d810b",
  1076 => x"80c9a80c",
  1077 => x"8454d008",
  1078 => x"708f2a70",
  1079 => x"81065151",
  1080 => x"5372f338",
  1081 => x"72d00ca0",
  1082 => x"f92dbff4",
  1083 => x"5186c52d",
  1084 => x"d008708f",
  1085 => x"2a708106",
  1086 => x"51515372",
  1087 => x"f338810b",
  1088 => x"d00cb153",
  1089 => x"805284d4",
  1090 => x"80c051a0",
  1091 => x"862d80c8",
  1092 => x"b408812e",
  1093 => x"93387282",
  1094 => x"2ebf38ff",
  1095 => x"135372e4",
  1096 => x"38ff1454",
  1097 => x"73ffaf38",
  1098 => x"a0f92d83",
  1099 => x"aa52849c",
  1100 => x"80c851a0",
  1101 => x"862d80c8",
  1102 => x"b408812e",
  1103 => x"09810693",
  1104 => x"389fb72d",
  1105 => x"80c8b408",
  1106 => x"83ffff06",
  1107 => x"537283aa",
  1108 => x"2e9f38a1",
  1109 => x"922da2ec",
  1110 => x"0480c080",
  1111 => x"5186c52d",
  1112 => x"8053a4c1",
  1113 => x"0480c098",
  1114 => x"5186c52d",
  1115 => x"8054a492",
  1116 => x"0481ff0b",
  1117 => x"d40cb154",
  1118 => x"a0f92d8f",
  1119 => x"cf538052",
  1120 => x"87fc80f7",
  1121 => x"51a0862d",
  1122 => x"80c8b408",
  1123 => x"5580c8b4",
  1124 => x"08812e09",
  1125 => x"81069c38",
  1126 => x"81ff0bd4",
  1127 => x"0c820a52",
  1128 => x"849c80e9",
  1129 => x"51a0862d",
  1130 => x"80c8b408",
  1131 => x"802e8d38",
  1132 => x"a0f92dff",
  1133 => x"135372c6",
  1134 => x"38a48504",
  1135 => x"81ff0bd4",
  1136 => x"0c80c8b4",
  1137 => x"085287fc",
  1138 => x"80fa51a0",
  1139 => x"862d80c8",
  1140 => x"b408b238",
  1141 => x"81ff0bd4",
  1142 => x"0cd40853",
  1143 => x"81ff0bd4",
  1144 => x"0c81ff0b",
  1145 => x"d40c81ff",
  1146 => x"0bd40c81",
  1147 => x"ff0bd40c",
  1148 => x"72862a70",
  1149 => x"81067656",
  1150 => x"51537296",
  1151 => x"3880c8b4",
  1152 => x"0854a492",
  1153 => x"0473822e",
  1154 => x"fedb38ff",
  1155 => x"145473fe",
  1156 => x"e7387380",
  1157 => x"c9a80c73",
  1158 => x"8b388152",
  1159 => x"87fc80d0",
  1160 => x"51a0862d",
  1161 => x"81ff0bd4",
  1162 => x"0cd00870",
  1163 => x"8f2a7081",
  1164 => x"06515153",
  1165 => x"72f33872",
  1166 => x"d00c81ff",
  1167 => x"0bd40c81",
  1168 => x"537280c8",
  1169 => x"b40c0294",
  1170 => x"050d0402",
  1171 => x"e8050d78",
  1172 => x"55805681",
  1173 => x"ff0bd40c",
  1174 => x"d008708f",
  1175 => x"2a708106",
  1176 => x"51515372",
  1177 => x"f3388281",
  1178 => x"0bd00c81",
  1179 => x"ff0bd40c",
  1180 => x"775287fc",
  1181 => x"80d151a0",
  1182 => x"862d80db",
  1183 => x"c6df5480",
  1184 => x"c8b40880",
  1185 => x"2e8b3880",
  1186 => x"c0b85186",
  1187 => x"c52da5e5",
  1188 => x"0481ff0b",
  1189 => x"d40cd408",
  1190 => x"7081ff06",
  1191 => x"51537281",
  1192 => x"fe2e0981",
  1193 => x"069e3880",
  1194 => x"ff539fb7",
  1195 => x"2d80c8b4",
  1196 => x"08757084",
  1197 => x"05570cff",
  1198 => x"13537280",
  1199 => x"25ec3881",
  1200 => x"56a5ca04",
  1201 => x"ff145473",
  1202 => x"c83881ff",
  1203 => x"0bd40c81",
  1204 => x"ff0bd40c",
  1205 => x"d008708f",
  1206 => x"2a708106",
  1207 => x"51515372",
  1208 => x"f33872d0",
  1209 => x"0c7580c8",
  1210 => x"b40c0298",
  1211 => x"050d0402",
  1212 => x"e8050d77",
  1213 => x"797b5855",
  1214 => x"55805372",
  1215 => x"7625a338",
  1216 => x"74708105",
  1217 => x"5680f52d",
  1218 => x"74708105",
  1219 => x"5680f52d",
  1220 => x"52527171",
  1221 => x"2e863881",
  1222 => x"51a6a404",
  1223 => x"811353a5",
  1224 => x"fb048051",
  1225 => x"7080c8b4",
  1226 => x"0c029805",
  1227 => x"0d0402ec",
  1228 => x"050d7655",
  1229 => x"74802e80",
  1230 => x"c2389a15",
  1231 => x"80e02d51",
  1232 => x"b4c32d80",
  1233 => x"c8b40880",
  1234 => x"c8b40880",
  1235 => x"cfdc0c80",
  1236 => x"c8b40854",
  1237 => x"5480cfb8",
  1238 => x"08802e9a",
  1239 => x"38941580",
  1240 => x"e02d51b4",
  1241 => x"c32d80c8",
  1242 => x"b408902b",
  1243 => x"83fff00a",
  1244 => x"06707507",
  1245 => x"51537280",
  1246 => x"cfdc0c80",
  1247 => x"cfdc0853",
  1248 => x"72802e9d",
  1249 => x"3880cfb0",
  1250 => x"08fe1471",
  1251 => x"2980cfc4",
  1252 => x"080580cf",
  1253 => x"e00c7084",
  1254 => x"2b80cfbc",
  1255 => x"0c54a7cf",
  1256 => x"0480cfc8",
  1257 => x"0880cfdc",
  1258 => x"0c80cfcc",
  1259 => x"0880cfe0",
  1260 => x"0c80cfb8",
  1261 => x"08802e8b",
  1262 => x"3880cfb0",
  1263 => x"08842b53",
  1264 => x"a7ca0480",
  1265 => x"cfd00884",
  1266 => x"2b537280",
  1267 => x"cfbc0c02",
  1268 => x"94050d04",
  1269 => x"02d8050d",
  1270 => x"800b80cf",
  1271 => x"b80c8454",
  1272 => x"a1ca2d80",
  1273 => x"c8b40880",
  1274 => x"2e973880",
  1275 => x"c9ac5280",
  1276 => x"51a4cb2d",
  1277 => x"80c8b408",
  1278 => x"802e8638",
  1279 => x"fe54a889",
  1280 => x"04ff1454",
  1281 => x"738024d8",
  1282 => x"38738d38",
  1283 => x"80c0c851",
  1284 => x"86c52d73",
  1285 => x"55adde04",
  1286 => x"8056810b",
  1287 => x"80cfe40c",
  1288 => x"885380c0",
  1289 => x"dc5280c9",
  1290 => x"e251a5ef",
  1291 => x"2d80c8b4",
  1292 => x"08762e09",
  1293 => x"81068938",
  1294 => x"80c8b408",
  1295 => x"80cfe40c",
  1296 => x"885380c0",
  1297 => x"e85280c9",
  1298 => x"fe51a5ef",
  1299 => x"2d80c8b4",
  1300 => x"08893880",
  1301 => x"c8b40880",
  1302 => x"cfe40c80",
  1303 => x"cfe40880",
  1304 => x"2e818138",
  1305 => x"80ccf20b",
  1306 => x"80f52d80",
  1307 => x"ccf30b80",
  1308 => x"f52d7198",
  1309 => x"2b71902b",
  1310 => x"0780ccf4",
  1311 => x"0b80f52d",
  1312 => x"70882b72",
  1313 => x"0780ccf5",
  1314 => x"0b80f52d",
  1315 => x"710780cd",
  1316 => x"aa0b80f5",
  1317 => x"2d80cdab",
  1318 => x"0b80f52d",
  1319 => x"71882b07",
  1320 => x"535f5452",
  1321 => x"5a565755",
  1322 => x"7381abaa",
  1323 => x"2e098106",
  1324 => x"8e387551",
  1325 => x"b4922d80",
  1326 => x"c8b40856",
  1327 => x"a9cd0473",
  1328 => x"82d4d52e",
  1329 => x"883880c0",
  1330 => x"f451aa99",
  1331 => x"0480c9ac",
  1332 => x"527551a4",
  1333 => x"cb2d80c8",
  1334 => x"b4085580",
  1335 => x"c8b40880",
  1336 => x"2e83fb38",
  1337 => x"885380c0",
  1338 => x"e85280c9",
  1339 => x"fe51a5ef",
  1340 => x"2d80c8b4",
  1341 => x"088a3881",
  1342 => x"0b80cfb8",
  1343 => x"0caa9f04",
  1344 => x"885380c0",
  1345 => x"dc5280c9",
  1346 => x"e251a5ef",
  1347 => x"2d80c8b4",
  1348 => x"08802e8b",
  1349 => x"3880c188",
  1350 => x"5186c52d",
  1351 => x"aafe0480",
  1352 => x"cdaa0b80",
  1353 => x"f52d5473",
  1354 => x"80d52e09",
  1355 => x"810680ce",
  1356 => x"3880cdab",
  1357 => x"0b80f52d",
  1358 => x"547381aa",
  1359 => x"2e098106",
  1360 => x"bd38800b",
  1361 => x"80c9ac0b",
  1362 => x"80f52d56",
  1363 => x"547481e9",
  1364 => x"2e833881",
  1365 => x"547481eb",
  1366 => x"2e8c3880",
  1367 => x"5573752e",
  1368 => x"09810682",
  1369 => x"f93880c9",
  1370 => x"b70b80f5",
  1371 => x"2d55748e",
  1372 => x"3880c9b8",
  1373 => x"0b80f52d",
  1374 => x"5473822e",
  1375 => x"86388055",
  1376 => x"adde0480",
  1377 => x"c9b90b80",
  1378 => x"f52d7080",
  1379 => x"cfb00cff",
  1380 => x"0580cfb4",
  1381 => x"0c80c9ba",
  1382 => x"0b80f52d",
  1383 => x"80c9bb0b",
  1384 => x"80f52d58",
  1385 => x"76057782",
  1386 => x"80290570",
  1387 => x"80cfc00c",
  1388 => x"80c9bc0b",
  1389 => x"80f52d70",
  1390 => x"80cfd40c",
  1391 => x"80cfb808",
  1392 => x"59575876",
  1393 => x"802e81b7",
  1394 => x"38885380",
  1395 => x"c0e85280",
  1396 => x"c9fe51a5",
  1397 => x"ef2d80c8",
  1398 => x"b4088282",
  1399 => x"3880cfb0",
  1400 => x"0870842b",
  1401 => x"80cfbc0c",
  1402 => x"7080cfd0",
  1403 => x"0c80c9d1",
  1404 => x"0b80f52d",
  1405 => x"80c9d00b",
  1406 => x"80f52d71",
  1407 => x"82802905",
  1408 => x"80c9d20b",
  1409 => x"80f52d70",
  1410 => x"84808029",
  1411 => x"1280c9d3",
  1412 => x"0b80f52d",
  1413 => x"7081800a",
  1414 => x"29127080",
  1415 => x"cfd80c80",
  1416 => x"cfd40871",
  1417 => x"2980cfc0",
  1418 => x"08057080",
  1419 => x"cfc40c80",
  1420 => x"c9d90b80",
  1421 => x"f52d80c9",
  1422 => x"d80b80f5",
  1423 => x"2d718280",
  1424 => x"290580c9",
  1425 => x"da0b80f5",
  1426 => x"2d708480",
  1427 => x"80291280",
  1428 => x"c9db0b80",
  1429 => x"f52d7098",
  1430 => x"2b81f00a",
  1431 => x"06720570",
  1432 => x"80cfc80c",
  1433 => x"fe117e29",
  1434 => x"770580cf",
  1435 => x"cc0c5259",
  1436 => x"5243545e",
  1437 => x"51525952",
  1438 => x"5d575957",
  1439 => x"add70480",
  1440 => x"c9be0b80",
  1441 => x"f52d80c9",
  1442 => x"bd0b80f5",
  1443 => x"2d718280",
  1444 => x"29057080",
  1445 => x"cfbc0c70",
  1446 => x"a02983ff",
  1447 => x"0570892a",
  1448 => x"7080cfd0",
  1449 => x"0c80c9c3",
  1450 => x"0b80f52d",
  1451 => x"80c9c20b",
  1452 => x"80f52d71",
  1453 => x"82802905",
  1454 => x"7080cfd8",
  1455 => x"0c7b7129",
  1456 => x"1e7080cf",
  1457 => x"cc0c7d80",
  1458 => x"cfc80c73",
  1459 => x"0580cfc4",
  1460 => x"0c555e51",
  1461 => x"51555580",
  1462 => x"51a6ae2d",
  1463 => x"81557480",
  1464 => x"c8b40c02",
  1465 => x"a8050d04",
  1466 => x"02ec050d",
  1467 => x"7670872c",
  1468 => x"7180ff06",
  1469 => x"55565480",
  1470 => x"cfb8088a",
  1471 => x"3873882c",
  1472 => x"7481ff06",
  1473 => x"545580c9",
  1474 => x"ac5280cf",
  1475 => x"c0081551",
  1476 => x"a4cb2d80",
  1477 => x"c8b40854",
  1478 => x"80c8b408",
  1479 => x"802eb838",
  1480 => x"80cfb808",
  1481 => x"802e9a38",
  1482 => x"72842980",
  1483 => x"c9ac0570",
  1484 => x"085253b4",
  1485 => x"922d80c8",
  1486 => x"b408f00a",
  1487 => x"0653aed5",
  1488 => x"04721080",
  1489 => x"c9ac0570",
  1490 => x"80e02d52",
  1491 => x"53b4c32d",
  1492 => x"80c8b408",
  1493 => x"53725473",
  1494 => x"80c8b40c",
  1495 => x"0294050d",
  1496 => x"0402e005",
  1497 => x"0d797084",
  1498 => x"2c80cfe0",
  1499 => x"0805718f",
  1500 => x"06525553",
  1501 => x"728a3880",
  1502 => x"c9ac5273",
  1503 => x"51a4cb2d",
  1504 => x"72a02980",
  1505 => x"c9ac0554",
  1506 => x"807480f5",
  1507 => x"2d565374",
  1508 => x"732e8338",
  1509 => x"81537481",
  1510 => x"e52e81f4",
  1511 => x"38817074",
  1512 => x"06545872",
  1513 => x"802e81e8",
  1514 => x"388b1480",
  1515 => x"f52d7083",
  1516 => x"2a790658",
  1517 => x"56769b38",
  1518 => x"80c6f808",
  1519 => x"53728938",
  1520 => x"7280cdac",
  1521 => x"0b81b72d",
  1522 => x"7680c6f8",
  1523 => x"0c7353b1",
  1524 => x"9204758f",
  1525 => x"2e098106",
  1526 => x"81b63874",
  1527 => x"9f068d29",
  1528 => x"80cd9f11",
  1529 => x"51538114",
  1530 => x"80f52d73",
  1531 => x"70810555",
  1532 => x"81b72d83",
  1533 => x"1480f52d",
  1534 => x"73708105",
  1535 => x"5581b72d",
  1536 => x"851480f5",
  1537 => x"2d737081",
  1538 => x"055581b7",
  1539 => x"2d871480",
  1540 => x"f52d7370",
  1541 => x"81055581",
  1542 => x"b72d8914",
  1543 => x"80f52d73",
  1544 => x"70810555",
  1545 => x"81b72d8e",
  1546 => x"1480f52d",
  1547 => x"73708105",
  1548 => x"5581b72d",
  1549 => x"901480f5",
  1550 => x"2d737081",
  1551 => x"055581b7",
  1552 => x"2d921480",
  1553 => x"f52d7370",
  1554 => x"81055581",
  1555 => x"b72d9414",
  1556 => x"80f52d73",
  1557 => x"70810555",
  1558 => x"81b72d96",
  1559 => x"1480f52d",
  1560 => x"73708105",
  1561 => x"5581b72d",
  1562 => x"981480f5",
  1563 => x"2d737081",
  1564 => x"055581b7",
  1565 => x"2d9c1480",
  1566 => x"f52d7370",
  1567 => x"81055581",
  1568 => x"b72d9e14",
  1569 => x"80f52d73",
  1570 => x"81b72d77",
  1571 => x"80c6f80c",
  1572 => x"80537280",
  1573 => x"c8b40c02",
  1574 => x"a0050d04",
  1575 => x"02cc050d",
  1576 => x"7e605e5a",
  1577 => x"800b80cf",
  1578 => x"dc0880cf",
  1579 => x"e008595c",
  1580 => x"56805880",
  1581 => x"cfbc0878",
  1582 => x"2e81b838",
  1583 => x"778f06a0",
  1584 => x"17575473",
  1585 => x"913880c9",
  1586 => x"ac527651",
  1587 => x"811757a4",
  1588 => x"cb2d80c9",
  1589 => x"ac568076",
  1590 => x"80f52d56",
  1591 => x"5474742e",
  1592 => x"83388154",
  1593 => x"7481e52e",
  1594 => x"80fd3881",
  1595 => x"70750655",
  1596 => x"5c73802e",
  1597 => x"80f1388b",
  1598 => x"1680f52d",
  1599 => x"98065978",
  1600 => x"80e5388b",
  1601 => x"537c5275",
  1602 => x"51a5ef2d",
  1603 => x"80c8b408",
  1604 => x"80d5389c",
  1605 => x"160851b4",
  1606 => x"922d80c8",
  1607 => x"b408841b",
  1608 => x"0c9a1680",
  1609 => x"e02d51b4",
  1610 => x"c32d80c8",
  1611 => x"b40880c8",
  1612 => x"b408881c",
  1613 => x"0c80c8b4",
  1614 => x"08555580",
  1615 => x"cfb80880",
  1616 => x"2e993894",
  1617 => x"1680e02d",
  1618 => x"51b4c32d",
  1619 => x"80c8b408",
  1620 => x"902b83ff",
  1621 => x"f00a0670",
  1622 => x"16515473",
  1623 => x"881b0c78",
  1624 => x"7a0c7b54",
  1625 => x"b3af0481",
  1626 => x"185880cf",
  1627 => x"bc087826",
  1628 => x"feca3880",
  1629 => x"cfb80880",
  1630 => x"2eb3387a",
  1631 => x"51ade82d",
  1632 => x"80c8b408",
  1633 => x"80c8b408",
  1634 => x"80ffffff",
  1635 => x"f806555b",
  1636 => x"7380ffff",
  1637 => x"fff82e95",
  1638 => x"3880c8b4",
  1639 => x"08fe0580",
  1640 => x"cfb00829",
  1641 => x"80cfc408",
  1642 => x"0557b1b1",
  1643 => x"04805473",
  1644 => x"80c8b40c",
  1645 => x"02b4050d",
  1646 => x"0402f405",
  1647 => x"0d747008",
  1648 => x"8105710c",
  1649 => x"700880cf",
  1650 => x"b4080653",
  1651 => x"53718f38",
  1652 => x"88130851",
  1653 => x"ade82d80",
  1654 => x"c8b40888",
  1655 => x"140c810b",
  1656 => x"80c8b40c",
  1657 => x"028c050d",
  1658 => x"0402f005",
  1659 => x"0d758811",
  1660 => x"08fe0580",
  1661 => x"cfb00829",
  1662 => x"80cfc408",
  1663 => x"11720880",
  1664 => x"cfb40806",
  1665 => x"05795553",
  1666 => x"5454a4cb",
  1667 => x"2d029005",
  1668 => x"0d0402f4",
  1669 => x"050d7470",
  1670 => x"882a83fe",
  1671 => x"80067072",
  1672 => x"982a0772",
  1673 => x"882b87fc",
  1674 => x"80800673",
  1675 => x"982b81f0",
  1676 => x"0a067173",
  1677 => x"070780c8",
  1678 => x"b40c5651",
  1679 => x"5351028c",
  1680 => x"050d0402",
  1681 => x"f8050d02",
  1682 => x"8e0580f5",
  1683 => x"2d74882b",
  1684 => x"077083ff",
  1685 => x"ff0680c8",
  1686 => x"b40c5102",
  1687 => x"88050d04",
  1688 => x"02f4050d",
  1689 => x"74767853",
  1690 => x"54528071",
  1691 => x"25973872",
  1692 => x"70810554",
  1693 => x"80f52d72",
  1694 => x"70810554",
  1695 => x"81b72dff",
  1696 => x"115170eb",
  1697 => x"38807281",
  1698 => x"b72d028c",
  1699 => x"050d0402",
  1700 => x"e8050d77",
  1701 => x"56807056",
  1702 => x"54737624",
  1703 => x"b63880cf",
  1704 => x"bc08742e",
  1705 => x"ae387351",
  1706 => x"aee12d80",
  1707 => x"c8b40880",
  1708 => x"c8b40809",
  1709 => x"81057080",
  1710 => x"c8b40807",
  1711 => x"9f2a7705",
  1712 => x"81175757",
  1713 => x"53537476",
  1714 => x"24893880",
  1715 => x"cfbc0874",
  1716 => x"26d43872",
  1717 => x"80c8b40c",
  1718 => x"0298050d",
  1719 => x"0402ec05",
  1720 => x"0d80c8b0",
  1721 => x"081751b5",
  1722 => x"8f2d80c8",
  1723 => x"b4085580",
  1724 => x"c8b40880",
  1725 => x"2ea2388b",
  1726 => x"5380c8b4",
  1727 => x"085280cd",
  1728 => x"ac51b4e0",
  1729 => x"2d80cfe8",
  1730 => x"08547380",
  1731 => x"2e8a3888",
  1732 => x"155280cd",
  1733 => x"ac51732d",
  1734 => x"0294050d",
  1735 => x"0402dc05",
  1736 => x"0d80705a",
  1737 => x"557480c8",
  1738 => x"b00825b4",
  1739 => x"3880cfbc",
  1740 => x"08752eac",
  1741 => x"387851ae",
  1742 => x"e12d80c8",
  1743 => x"b4080981",
  1744 => x"057080c8",
  1745 => x"b408079f",
  1746 => x"2a760581",
  1747 => x"1b5b5654",
  1748 => x"7480c8b0",
  1749 => x"08258938",
  1750 => x"80cfbc08",
  1751 => x"7926d638",
  1752 => x"80557880",
  1753 => x"cfbc0827",
  1754 => x"81db3878",
  1755 => x"51aee12d",
  1756 => x"80c8b408",
  1757 => x"802e81ad",
  1758 => x"3880c8b4",
  1759 => x"088b0580",
  1760 => x"f52d7084",
  1761 => x"2a708106",
  1762 => x"77107884",
  1763 => x"2b80cdac",
  1764 => x"0b80f52d",
  1765 => x"5c5c5351",
  1766 => x"55567380",
  1767 => x"2e80cb38",
  1768 => x"7416822b",
  1769 => x"b8e90b80",
  1770 => x"c784120c",
  1771 => x"54777531",
  1772 => x"1080cfec",
  1773 => x"11555690",
  1774 => x"74708105",
  1775 => x"5681b72d",
  1776 => x"a07481b7",
  1777 => x"2d7681ff",
  1778 => x"06811658",
  1779 => x"5473802e",
  1780 => x"8a389c53",
  1781 => x"80cdac52",
  1782 => x"b7e2048b",
  1783 => x"5380c8b4",
  1784 => x"085280cf",
  1785 => x"ee1651b8",
  1786 => x"9d047416",
  1787 => x"822bb5dd",
  1788 => x"0b80c784",
  1789 => x"120c5476",
  1790 => x"81ff0681",
  1791 => x"16585473",
  1792 => x"802e8a38",
  1793 => x"9c5380cd",
  1794 => x"ac52b894",
  1795 => x"048b5380",
  1796 => x"c8b40852",
  1797 => x"77753110",
  1798 => x"80cfec05",
  1799 => x"517655b4",
  1800 => x"e02db8ba",
  1801 => x"04749029",
  1802 => x"75317010",
  1803 => x"80cfec05",
  1804 => x"515480c8",
  1805 => x"b4087481",
  1806 => x"b72d8119",
  1807 => x"59748b24",
  1808 => x"a338b6e2",
  1809 => x"04749029",
  1810 => x"75317010",
  1811 => x"80cfec05",
  1812 => x"8c773157",
  1813 => x"51548074",
  1814 => x"81b72d9e",
  1815 => x"14ff1656",
  1816 => x"5474f338",
  1817 => x"02a4050d",
  1818 => x"0402fc05",
  1819 => x"0d80c8b0",
  1820 => x"081351b5",
  1821 => x"8f2d80c8",
  1822 => x"b408802e",
  1823 => x"893880c8",
  1824 => x"b40851a6",
  1825 => x"ae2d800b",
  1826 => x"80c8b00c",
  1827 => x"b69d2d91",
  1828 => x"832d0284",
  1829 => x"050d0402",
  1830 => x"fc050d72",
  1831 => x"5170fd2e",
  1832 => x"b03870fd",
  1833 => x"248a3870",
  1834 => x"fc2e80cc",
  1835 => x"38ba8204",
  1836 => x"70fe2eb7",
  1837 => x"3870ff2e",
  1838 => x"09810680",
  1839 => x"c53880c8",
  1840 => x"b0085170",
  1841 => x"802ebb38",
  1842 => x"ff1180c8",
  1843 => x"b00cba82",
  1844 => x"0480c8b0",
  1845 => x"08f40570",
  1846 => x"80c8b00c",
  1847 => x"51708025",
  1848 => x"a138800b",
  1849 => x"80c8b00c",
  1850 => x"ba820480",
  1851 => x"c8b00881",
  1852 => x"0580c8b0",
  1853 => x"0cba8204",
  1854 => x"80c8b008",
  1855 => x"8c0580c8",
  1856 => x"b00cb69d",
  1857 => x"2d91832d",
  1858 => x"0284050d",
  1859 => x"0402fc05",
  1860 => x"0d800b80",
  1861 => x"c8b00cb6",
  1862 => x"9d2d8ff1",
  1863 => x"2d80c8b4",
  1864 => x"0880c8a0",
  1865 => x"0c80c6fc",
  1866 => x"5192a62d",
  1867 => x"0284050d",
  1868 => x"047180cf",
  1869 => x"e80c0400",
  1870 => x"00ffffff",
  1871 => x"ff00ffff",
  1872 => x"ffff00ff",
  1873 => x"ffffff00",
  1874 => x"20204368",
  1875 => x"69702d38",
  1876 => x"3a202020",
  1877 => x"20202020",
  1878 => x"50532f32",
  1879 => x"3a000000",
  1880 => x"20203120",
  1881 => x"32203320",
  1882 => x"43202020",
  1883 => x"20202020",
  1884 => x"31203220",
  1885 => x"33203400",
  1886 => x"20203420",
  1887 => x"35203620",
  1888 => x"44202020",
  1889 => x"20202020",
  1890 => x"51205720",
  1891 => x"45205200",
  1892 => x"20203720",
  1893 => x"38203920",
  1894 => x"45202020",
  1895 => x"20202020",
  1896 => x"41205320",
  1897 => x"44204600",
  1898 => x"20204120",
  1899 => x"30204220",
  1900 => x"46202020",
  1901 => x"20202020",
  1902 => x"5a205820",
  1903 => x"43205600",
  1904 => x"3d3d3d20",
  1905 => x"43484950",
  1906 => x"2d382066",
  1907 => x"6f72205a",
  1908 => x"58444f53",
  1909 => x"203d3d3d",
  1910 => x"00000000",
  1911 => x"52657365",
  1912 => x"74000000",
  1913 => x"4c6f6164",
  1914 => x"20526f6d",
  1915 => x"20282e62",
  1916 => x"696e2c20",
  1917 => x"2e636838",
  1918 => x"29201000",
  1919 => x"536f756e",
  1920 => x"64206f6e",
  1921 => x"2f6f6666",
  1922 => x"00000000",
  1923 => x"4b657962",
  1924 => x"6f617264",
  1925 => x"2048656c",
  1926 => x"70000000",
  1927 => x"45786974",
  1928 => x"00000000",
  1929 => x"436c6f63",
  1930 => x"6b205370",
  1931 => x"6565643a",
  1932 => x"20317800",
  1933 => x"436c6f63",
  1934 => x"6b205370",
  1935 => x"6565643a",
  1936 => x"20327800",
  1937 => x"436c6f63",
  1938 => x"6b205370",
  1939 => x"6565643a",
  1940 => x"20337800",
  1941 => x"436c6f63",
  1942 => x"6b205370",
  1943 => x"6565643a",
  1944 => x"20347800",
  1945 => x"3d3d3d20",
  1946 => x"43484950",
  1947 => x"2d382066",
  1948 => x"6f72205a",
  1949 => x"58554e4f",
  1950 => x"203d3d3d",
  1951 => x"00000000",
  1952 => x"524f4d20",
  1953 => x"6c6f6164",
  1954 => x"696e6720",
  1955 => x"6661696c",
  1956 => x"65640000",
  1957 => x"4f4b0000",
  1958 => x"3d3d3d20",
  1959 => x"43484950",
  1960 => x"2d38204b",
  1961 => x"6579626f",
  1962 => x"61726420",
  1963 => x"48454c50",
  1964 => x"203d3d3d",
  1965 => x"00000000",
  1966 => x"3d3d3d3d",
  1967 => x"3d3d3d3d",
  1968 => x"3d3d3d3d",
  1969 => x"3d3d3d3d",
  1970 => x"3d3d3d3d",
  1971 => x"3d3d3d3d",
  1972 => x"3d3d3d3d",
  1973 => x"00000000",
  1974 => x"43686970",
  1975 => x"2d382068",
  1976 => x"61732061",
  1977 => x"20686578",
  1978 => x"206b6579",
  1979 => x"7061642e",
  1980 => x"00000000",
  1981 => x"54686520",
  1982 => x"6d617070",
  1983 => x"696e6720",
  1984 => x"746f2050",
  1985 => x"43206b65",
  1986 => x"79626f61",
  1987 => x"72640000",
  1988 => x"69732066",
  1989 => x"6f6c6c6f",
  1990 => x"77696e67",
  1991 => x"2e000000",
  1992 => x"3d3d3d20",
  1993 => x"43484950",
  1994 => x"2d382043",
  1995 => x"6f726520",
  1996 => x"43726564",
  1997 => x"69747320",
  1998 => x"3d3d3d00",
  1999 => x"43686970",
  2000 => x"2d382063",
  2001 => x"6f726520",
  2002 => x"666f7220",
  2003 => x"5a58554e",
  2004 => x"4f2c2041",
  2005 => x"454f4e2c",
  2006 => x"00000000",
  2007 => x"5a58444f",
  2008 => x"5320616e",
  2009 => x"64205a58",
  2010 => x"444f532b",
  2011 => x"20626f61",
  2012 => x"7264732e",
  2013 => x"00000000",
  2014 => x"4f726967",
  2015 => x"696e616c",
  2016 => x"20636f72",
  2017 => x"65206279",
  2018 => x"3a000000",
  2019 => x"202d2043",
  2020 => x"61727374",
  2021 => x"656e2045",
  2022 => x"6c746f6e",
  2023 => x"20536f72",
  2024 => x"656e7365",
  2025 => x"6e200000",
  2026 => x"506f7274",
  2027 => x"206d6164",
  2028 => x"65206279",
  2029 => x"3a000000",
  2030 => x"202d2041",
  2031 => x"7a65736d",
  2032 => x"626f6700",
  2033 => x"202d2041",
  2034 => x"766c6978",
  2035 => x"41000000",
  2036 => x"496e6974",
  2037 => x"69616c69",
  2038 => x"7a696e67",
  2039 => x"20534420",
  2040 => x"63617264",
  2041 => x"0a000000",
  2042 => x"16200000",
  2043 => x"14200000",
  2044 => x"15200000",
  2045 => x"53442069",
  2046 => x"6e69742e",
  2047 => x"2e2e0a00",
  2048 => x"53442063",
  2049 => x"61726420",
  2050 => x"72657365",
  2051 => x"74206661",
  2052 => x"696c6564",
  2053 => x"210a0000",
  2054 => x"53444843",
  2055 => x"20657272",
  2056 => x"6f72210a",
  2057 => x"00000000",
  2058 => x"57726974",
  2059 => x"65206661",
  2060 => x"696c6564",
  2061 => x"0a000000",
  2062 => x"52656164",
  2063 => x"20666169",
  2064 => x"6c65640a",
  2065 => x"00000000",
  2066 => x"43617264",
  2067 => x"20696e69",
  2068 => x"74206661",
  2069 => x"696c6564",
  2070 => x"0a000000",
  2071 => x"46415431",
  2072 => x"36202020",
  2073 => x"00000000",
  2074 => x"46415433",
  2075 => x"32202020",
  2076 => x"00000000",
  2077 => x"4e6f2070",
  2078 => x"61727469",
  2079 => x"74696f6e",
  2080 => x"20736967",
  2081 => x"0a000000",
  2082 => x"42616420",
  2083 => x"70617274",
  2084 => x"0a000000",
  2085 => x"4261636b",
  2086 => x"00000000",
  2087 => x"00000002",
  2088 => x"00000000",
  2089 => x"00000002",
  2090 => x"00001dc0",
  2091 => x"000003ab",
  2092 => x"00000002",
  2093 => x"00001ebc",
  2094 => x"000003ab",
  2095 => x"00000002",
  2096 => x"00001ddc",
  2097 => x"0000037f",
  2098 => x"00000003",
  2099 => x"00002110",
  2100 => x"00000004",
  2101 => x"00000002",
  2102 => x"00001de4",
  2103 => x"00001d0d",
  2104 => x"00000001",
  2105 => x"00001dfc",
  2106 => x"00000000",
  2107 => x"00000002",
  2108 => x"00001e0c",
  2109 => x"000003c6",
  2110 => x"00000002",
  2111 => x"00001e1c",
  2112 => x"0000080e",
  2113 => x"00000000",
  2114 => x"00000000",
  2115 => x"00000000",
  2116 => x"00001e24",
  2117 => x"00001e34",
  2118 => x"00001e44",
  2119 => x"00001e54",
  2120 => x"00000002",
  2121 => x"00001e64",
  2122 => x"000003ab",
  2123 => x"00000002",
  2124 => x"00001ebc",
  2125 => x"000003ab",
  2126 => x"00000002",
  2127 => x"00001ddc",
  2128 => x"0000037f",
  2129 => x"00000003",
  2130 => x"00002110",
  2131 => x"00000004",
  2132 => x"00000002",
  2133 => x"00001de4",
  2134 => x"00001d0d",
  2135 => x"00000001",
  2136 => x"00001dfc",
  2137 => x"00000000",
  2138 => x"00000002",
  2139 => x"00001e0c",
  2140 => x"000003c6",
  2141 => x"00000002",
  2142 => x"00001e1c",
  2143 => x"0000080e",
  2144 => x"00000000",
  2145 => x"00000000",
  2146 => x"00000000",
  2147 => x"00000004",
  2148 => x"00001e80",
  2149 => x"0000218c",
  2150 => x"00000004",
  2151 => x"00001e94",
  2152 => x"00002460",
  2153 => x"00000000",
  2154 => x"00000000",
  2155 => x"00000000",
  2156 => x"00000002",
  2157 => x"00001e98",
  2158 => x"000003aa",
  2159 => x"00000002",
  2160 => x"00001eb8",
  2161 => x"000003aa",
  2162 => x"00000002",
  2163 => x"00001ed8",
  2164 => x"000003aa",
  2165 => x"00000002",
  2166 => x"00001ef4",
  2167 => x"000003aa",
  2168 => x"00000002",
  2169 => x"00001f10",
  2170 => x"000003aa",
  2171 => x"00000002",
  2172 => x"00002024",
  2173 => x"000003aa",
  2174 => x"00000002",
  2175 => x"00001d48",
  2176 => x"000003aa",
  2177 => x"00000002",
  2178 => x"00001d60",
  2179 => x"000003aa",
  2180 => x"00000002",
  2181 => x"00001d78",
  2182 => x"000003aa",
  2183 => x"00000002",
  2184 => x"00001d90",
  2185 => x"000003aa",
  2186 => x"00000002",
  2187 => x"00001da8",
  2188 => x"000003aa",
  2189 => x"00000002",
  2190 => x"00002024",
  2191 => x"000003aa",
  2192 => x"00000004",
  2193 => x"00001e94",
  2194 => x"00002460",
  2195 => x"00000000",
  2196 => x"00000000",
  2197 => x"00000000",
  2198 => x"00000002",
  2199 => x"00001f20",
  2200 => x"000003aa",
  2201 => x"00000002",
  2202 => x"00001eb8",
  2203 => x"000003aa",
  2204 => x"00000002",
  2205 => x"00001f3c",
  2206 => x"000003aa",
  2207 => x"00000002",
  2208 => x"00001f5c",
  2209 => x"000003aa",
  2210 => x"00000002",
  2211 => x"00002024",
  2212 => x"000003aa",
  2213 => x"00000002",
  2214 => x"00001f78",
  2215 => x"000003aa",
  2216 => x"00000002",
  2217 => x"00001f8c",
  2218 => x"000003aa",
  2219 => x"00000002",
  2220 => x"00002024",
  2221 => x"000003aa",
  2222 => x"00000002",
  2223 => x"00001fa8",
  2224 => x"000003aa",
  2225 => x"00000002",
  2226 => x"00001fb8",
  2227 => x"000003aa",
  2228 => x"00000002",
  2229 => x"00001fc4",
  2230 => x"000003aa",
  2231 => x"00000002",
  2232 => x"00002024",
  2233 => x"000003aa",
  2234 => x"00000004",
  2235 => x"00001e94",
  2236 => x"00002460",
  2237 => x"00000000",
  2238 => x"00000000",
  2239 => x"00000000",
  2240 => x"00000000",
  2241 => x"00000000",
  2242 => x"00000000",
  2243 => x"00000000",
  2244 => x"00000000",
  2245 => x"00000000",
  2246 => x"00000000",
  2247 => x"00000000",
  2248 => x"00000000",
  2249 => x"00000000",
  2250 => x"00000000",
  2251 => x"00000000",
  2252 => x"00000000",
  2253 => x"00000000",
  2254 => x"00000000",
  2255 => x"00000000",
  2256 => x"00000000",
  2257 => x"00000000",
  2258 => x"00000006",
  2259 => x"00000043",
  2260 => x"00000042",
  2261 => x"0000003b",
  2262 => x"0000004b",
  2263 => x"00000033",
  2264 => x"0000001d",
  2265 => x"0000001b",
  2266 => x"0000001c",
  2267 => x"00000023",
  2268 => x"0000002b",
  2269 => x"00000000",
  2270 => x"00000000",
  2271 => x"00000002",
  2272 => x"000027ec",
  2273 => x"00001add",
  2274 => x"00000002",
  2275 => x"0000280a",
  2276 => x"00001add",
  2277 => x"00000002",
  2278 => x"00002828",
  2279 => x"00001add",
  2280 => x"00000002",
  2281 => x"00002846",
  2282 => x"00001add",
  2283 => x"00000002",
  2284 => x"00002864",
  2285 => x"00001add",
  2286 => x"00000002",
  2287 => x"00002882",
  2288 => x"00001add",
  2289 => x"00000002",
  2290 => x"000028a0",
  2291 => x"00001add",
  2292 => x"00000002",
  2293 => x"000028be",
  2294 => x"00001add",
  2295 => x"00000002",
  2296 => x"000028dc",
  2297 => x"00001add",
  2298 => x"00000002",
  2299 => x"000028fa",
  2300 => x"00001add",
  2301 => x"00000002",
  2302 => x"00002918",
  2303 => x"00001add",
  2304 => x"00000002",
  2305 => x"00002936",
  2306 => x"00001add",
  2307 => x"00000002",
  2308 => x"00002954",
  2309 => x"00001add",
  2310 => x"00000004",
  2311 => x"00002094",
  2312 => x"00000000",
  2313 => x"00000000",
  2314 => x"00000000",
  2315 => x"00001c97",
  2316 => x"00000000",
	others => x"00000000"
);

begin

process (clk)
begin
	if (clk'event and clk = '1') then
		if (from_zpu.memAWriteEnable = '1') and (from_zpu.memBWriteEnable = '1') and (from_zpu.memAAddr=from_zpu.memBAddr) and (from_zpu.memAWrite/=from_zpu.memBWrite) then
			report "write collision" severity failure;
		end if;
	
		if (from_zpu.memAWriteEnable = '1') then
			ram(to_integer(unsigned(from_zpu.memAAddr(maxAddrBitBRAM downto 2)))) := from_zpu.memAWrite;
			to_zpu.memARead <= from_zpu.memAWrite;
		else
			to_zpu.memARead <= ram(to_integer(unsigned(from_zpu.memAAddr(maxAddrBitBRAM downto 2))));
		end if;
	end if;
end process;

process (clk)
begin
	if (clk'event and clk = '1') then
		if (from_zpu.memBWriteEnable = '1') then
			ram(to_integer(unsigned(from_zpu.memBAddr(maxAddrBitBRAM downto 2)))) := from_zpu.memBWrite;
			to_zpu.memBRead <= from_zpu.memBWrite;
		else
			to_zpu.memBRead <= ram(to_integer(unsigned(from_zpu.memBAddr(maxAddrBitBRAM downto 2))));
		end if;
	end if;
end process;


end arch;

