-- ZPU
--
-- Copyright 2004-2008 oharboe - �yvind Harboe - oyvind.harboe@zylin.com
-- Modified by Alastair M. Robinson for the ZPUFlex project.
--
-- The FreeBSD license
-- 
-- Redistribution and use in source and binary forms, with or without
-- modification, are permitted provided that the following conditions
-- are met:
-- 
-- 1. Redistributions of source code must retain the above copyright
--    notice, this list of conditions and the following disclaimer.
-- 2. Redistributions in binary form must reproduce the above
--    copyright notice, this list of conditions and the following
--    disclaimer in the documentation and/or other materials
--    provided with the distribution.
-- 
-- THIS SOFTWARE IS PROVIDED BY THE ZPU PROJECT ``AS IS'' AND ANY
-- EXPRESS OR IMPLIED WARRANTIES, INCLUDING, BUT NOT LIMITED TO,
-- THE IMPLIED WARRANTIES OF MERCHANTABILITY AND FITNESS FOR A
-- PARTICULAR PURPOSE ARE DISCLAIMED. IN NO EVENT SHALL THE
-- ZPU PROJECT OR CONTRIBUTORS BE LIABLE FOR ANY DIRECT,
-- INDIRECT, INCIDENTAL, SPECIAL, EXEMPLARY, OR CONSEQUENTIAL DAMAGES
-- (INCLUDING, BUT NOT LIMITED TO, PROCUREMENT OF SUBSTITUTE GOODS
-- OR SERVICES; LOSS OF USE, DATA, OR PROFITS; OR BUSINESS INTERRUPTION)
-- HOWEVER CAUSED AND ON ANY THEORY OF LIABILITY, WHETHER IN CONTRACT,
-- STRICT LIABILITY, OR TORT (INCLUDING NEGLIGENCE OR OTHERWISE)
-- ARISING IN ANY WAY OUT OF THE USE OF THIS SOFTWARE, EVEN IF
-- ADVISED OF THE POSSIBILITY OF SUCH DAMAGE.
-- 
-- The views and conclusions contained in the software and documentation
-- are those of the authors and should not be interpreted as representing
-- official policies, either expressed or implied, of the ZPU Project.

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;


library work;
use work.zpupkg.all;

entity CtrlROM_ROM is
generic
	(
		maxAddrBitBRAM : integer := maxAddrBitBRAMLimit -- Specify your actual ROM size to save LEs and unnecessary block RAM usage.
	);
port (
	clk : in std_logic;
	areset : in std_logic := '0';
	from_zpu : in ZPU_ToROM;
	to_zpu : out ZPU_FromROM
);
end CtrlROM_ROM;

architecture arch of CtrlROM_ROM is

type ram_type is array(natural range 0 to ((2**(maxAddrBitBRAM+1))/4)-1) of std_logic_vector(wordSize-1 downto 0);

shared variable ram : ram_type :=
(
     0 => x"0b0b0b0b",
     1 => x"8c0b0b0b",
     2 => x"0b81e004",
     3 => x"0b0b0b0b",
     4 => x"8c04ff0d",
     5 => x"80040400",
     6 => x"00000016",
     7 => x"00000000",
     8 => x"0b0b0bab",
     9 => x"ec080b0b",
    10 => x"0babf008",
    11 => x"0b0b0bab",
    12 => x"f4080b0b",
    13 => x"0b0b9808",
    14 => x"2d0b0b0b",
    15 => x"abf40c0b",
    16 => x"0b0babf0",
    17 => x"0c0b0b0b",
    18 => x"abec0c04",
    19 => x"00000000",
    20 => x"00000000",
    21 => x"00000000",
    22 => x"00000000",
    23 => x"00000000",
    24 => x"71fd0608",
    25 => x"72830609",
    26 => x"81058205",
    27 => x"832b2a83",
    28 => x"ffff0652",
    29 => x"0471fc06",
    30 => x"08728306",
    31 => x"09810583",
    32 => x"05101010",
    33 => x"2a81ff06",
    34 => x"520471fd",
    35 => x"060883ff",
    36 => x"ff738306",
    37 => x"09810582",
    38 => x"05832b2b",
    39 => x"09067383",
    40 => x"ffff0673",
    41 => x"83060981",
    42 => x"05820583",
    43 => x"2b0b2b07",
    44 => x"72fc060c",
    45 => x"51510471",
    46 => x"fc06080b",
    47 => x"0b0ba688",
    48 => x"73830610",
    49 => x"10050806",
    50 => x"7381ff06",
    51 => x"73830609",
    52 => x"81058305",
    53 => x"1010102b",
    54 => x"0772fc06",
    55 => x"0c515104",
    56 => x"abec70b1",
    57 => x"88278b38",
    58 => x"80717084",
    59 => x"05530c81",
    60 => x"e2048c51",
    61 => x"85e80402",
    62 => x"fc050df8",
    63 => x"80518f0b",
    64 => x"abfc0c9f",
    65 => x"0bac800c",
    66 => x"a0717081",
    67 => x"055334ac",
    68 => x"8008ff05",
    69 => x"ac800cac",
    70 => x"80088025",
    71 => x"eb38abfc",
    72 => x"08ff05ab",
    73 => x"fc0cabfc",
    74 => x"088025d7",
    75 => x"38800bac",
    76 => x"800c800b",
    77 => x"abfc0c02",
    78 => x"84050d04",
    79 => x"02f0050d",
    80 => x"f88053f8",
    81 => x"a05483bf",
    82 => x"52737081",
    83 => x"05553351",
    84 => x"70737081",
    85 => x"055534ff",
    86 => x"12527180",
    87 => x"25eb38fb",
    88 => x"c0539f52",
    89 => x"a0737081",
    90 => x"055534ff",
    91 => x"12527180",
    92 => x"25f23802",
    93 => x"90050d04",
    94 => x"02f4050d",
    95 => x"74538e0b",
    96 => x"abfc0825",
    97 => x"8f3882bc",
    98 => x"2dabfc08",
    99 => x"ff05abfc",
   100 => x"0c82fe04",
   101 => x"abfc08ac",
   102 => x"80085351",
   103 => x"728a2e09",
   104 => x"8106b738",
   105 => x"7151719f",
   106 => x"24a038ab",
   107 => x"fc08a029",
   108 => x"11f88011",
   109 => x"5151a071",
   110 => x"34ac8008",
   111 => x"8105ac80",
   112 => x"0cac8008",
   113 => x"519f7125",
   114 => x"e238800b",
   115 => x"ac800cab",
   116 => x"fc088105",
   117 => x"abfc0c83",
   118 => x"ee0470a0",
   119 => x"2912f880",
   120 => x"11515172",
   121 => x"7134ac80",
   122 => x"088105ac",
   123 => x"800cac80",
   124 => x"08a02e09",
   125 => x"81068e38",
   126 => x"800bac80",
   127 => x"0cabfc08",
   128 => x"8105abfc",
   129 => x"0c028c05",
   130 => x"0d0402ec",
   131 => x"050d800b",
   132 => x"ac840cf6",
   133 => x"8c08f690",
   134 => x"0871882c",
   135 => x"565481ff",
   136 => x"06527372",
   137 => x"25883871",
   138 => x"54820bac",
   139 => x"840c7288",
   140 => x"2c7381ff",
   141 => x"06545574",
   142 => x"73258b38",
   143 => x"72ac8408",
   144 => x"8407ac84",
   145 => x"0c557384",
   146 => x"2b86a071",
   147 => x"25827131",
   148 => x"700b0b0b",
   149 => x"a9c00c81",
   150 => x"712bff05",
   151 => x"f6880cfc",
   152 => x"08fefe14",
   153 => x"ff132c79",
   154 => x"8829ff94",
   155 => x"0570812c",
   156 => x"ac840852",
   157 => x"59535155",
   158 => x"51525476",
   159 => x"802e8538",
   160 => x"70810751",
   161 => x"70f6940c",
   162 => x"71098105",
   163 => x"f6800c72",
   164 => x"098105f6",
   165 => x"840c0294",
   166 => x"050d0402",
   167 => x"f4050d74",
   168 => x"53727081",
   169 => x"055480f5",
   170 => x"2d527180",
   171 => x"2e893871",
   172 => x"5182f82d",
   173 => x"85a10481",
   174 => x"0babec0c",
   175 => x"028c050d",
   176 => x"0402fc05",
   177 => x"0d818080",
   178 => x"51c01151",
   179 => x"70fb3802",
   180 => x"84050d04",
   181 => x"02fc050d",
   182 => x"ec518371",
   183 => x"0c85c12d",
   184 => x"82710c02",
   185 => x"84050d04",
   186 => x"02f0050d",
   187 => x"805185d4",
   188 => x"2d840bec",
   189 => x"0c8ba32d",
   190 => x"87ea2d81",
   191 => x"f72d8352",
   192 => x"8b882d81",
   193 => x"51848a2d",
   194 => x"ff125271",
   195 => x"8025f138",
   196 => x"840bec0c",
   197 => x"a7fc5185",
   198 => x"9b2d9ff7",
   199 => x"2dabec08",
   200 => x"802e81b1",
   201 => x"389f0bab",
   202 => x"bc0c9f0b",
   203 => x"fc0ca9c4",
   204 => x"518dee2d",
   205 => x"8bd22d8b",
   206 => x"e52d87f6",
   207 => x"2d8dfe2d",
   208 => x"aaac0b80",
   209 => x"f52d7087",
   210 => x"2babbc08",
   211 => x"70810653",
   212 => x"56545271",
   213 => x"802e8538",
   214 => x"72810753",
   215 => x"73812a70",
   216 => x"81065152",
   217 => x"71802e85",
   218 => x"38728207",
   219 => x"5373822a",
   220 => x"70810651",
   221 => x"5271802e",
   222 => x"85387284",
   223 => x"07537383",
   224 => x"2a708106",
   225 => x"51527180",
   226 => x"2e853872",
   227 => x"88075373",
   228 => x"842a7081",
   229 => x"06515271",
   230 => x"802e8538",
   231 => x"72900753",
   232 => x"73852a70",
   233 => x"81065152",
   234 => x"71802e85",
   235 => x"3872a007",
   236 => x"5373862a",
   237 => x"70810651",
   238 => x"5271802e",
   239 => x"86387280",
   240 => x"c0075372",
   241 => x"fc0c8652",
   242 => x"abec0883",
   243 => x"38845271",
   244 => x"ec0c86ba",
   245 => x"04800bab",
   246 => x"ec0c0290",
   247 => x"050d0471",
   248 => x"980c04ff",
   249 => x"b008abec",
   250 => x"0c04810b",
   251 => x"ffb00c04",
   252 => x"800bffb0",
   253 => x"0c0402f4",
   254 => x"050d88f8",
   255 => x"04abec08",
   256 => x"81f02e09",
   257 => x"81068938",
   258 => x"810babb4",
   259 => x"0c88f804",
   260 => x"abec0881",
   261 => x"e02e0981",
   262 => x"06893881",
   263 => x"0babb80c",
   264 => x"88f804ab",
   265 => x"ec0852ab",
   266 => x"b808802e",
   267 => x"8838abec",
   268 => x"08818005",
   269 => x"5271842c",
   270 => x"728f0653",
   271 => x"53abb408",
   272 => x"802e9938",
   273 => x"728429aa",
   274 => x"f4057213",
   275 => x"81712b70",
   276 => x"09730806",
   277 => x"730c5153",
   278 => x"5388ee04",
   279 => x"728429aa",
   280 => x"f4057213",
   281 => x"83712b72",
   282 => x"0807720c",
   283 => x"5353800b",
   284 => x"abb80c80",
   285 => x"0babb40c",
   286 => x"ac885189",
   287 => x"f92dabec",
   288 => x"08ff24fe",
   289 => x"f838800b",
   290 => x"abec0c02",
   291 => x"8c050d04",
   292 => x"02f8050d",
   293 => x"aaf4528f",
   294 => x"51807270",
   295 => x"8405540c",
   296 => x"ff115170",
   297 => x"8025f238",
   298 => x"0288050d",
   299 => x"0402f005",
   300 => x"0d755187",
   301 => x"f02d7082",
   302 => x"2cfc06aa",
   303 => x"f4117210",
   304 => x"9e067108",
   305 => x"70722a70",
   306 => x"83068274",
   307 => x"2b700974",
   308 => x"06760c54",
   309 => x"51565753",
   310 => x"515387ea",
   311 => x"2d71abec",
   312 => x"0c029005",
   313 => x"0d0402fc",
   314 => x"050d7251",
   315 => x"80710c80",
   316 => x"0b84120c",
   317 => x"0284050d",
   318 => x"0402f005",
   319 => x"0d757008",
   320 => x"84120853",
   321 => x"5353ff54",
   322 => x"71712ea8",
   323 => x"3887f02d",
   324 => x"84130870",
   325 => x"84291488",
   326 => x"11700870",
   327 => x"81ff0684",
   328 => x"18088111",
   329 => x"8706841a",
   330 => x"0c535155",
   331 => x"51515187",
   332 => x"ea2d7154",
   333 => x"73abec0c",
   334 => x"0290050d",
   335 => x"0402f405",
   336 => x"0d87f02d",
   337 => x"e008708b",
   338 => x"2a708106",
   339 => x"51525370",
   340 => x"802e9d38",
   341 => x"ac880870",
   342 => x"8429ac90",
   343 => x"057481ff",
   344 => x"06710c51",
   345 => x"51ac8808",
   346 => x"81118706",
   347 => x"ac880c51",
   348 => x"728c2cbf",
   349 => x"06acb00c",
   350 => x"800bacb4",
   351 => x"0c87e32d",
   352 => x"87ea2d02",
   353 => x"8c050d04",
   354 => x"02fc050d",
   355 => x"87f02d81",
   356 => x"0bacb40c",
   357 => x"87ea2dac",
   358 => x"b4085170",
   359 => x"fa380284",
   360 => x"050d0402",
   361 => x"fc050dac",
   362 => x"885189e6",
   363 => x"2d89902d",
   364 => x"8abd5187",
   365 => x"df2d0284",
   366 => x"050d0402",
   367 => x"fc050d8f",
   368 => x"cf5185c1",
   369 => x"2dff1151",
   370 => x"708025f6",
   371 => x"38028405",
   372 => x"0d0402fc",
   373 => x"050d810b",
   374 => x"abe80c81",
   375 => x"51848a2d",
   376 => x"0284050d",
   377 => x"0402fc05",
   378 => x"0d8bef04",
   379 => x"87f62d80",
   380 => x"f65189ad",
   381 => x"2dabec08",
   382 => x"f33880da",
   383 => x"5189ad2d",
   384 => x"abec08e8",
   385 => x"38abe408",
   386 => x"5189ad2d",
   387 => x"abec08dc",
   388 => x"38abec08",
   389 => x"abe80cab",
   390 => x"ec085184",
   391 => x"8a2d0284",
   392 => x"050d0402",
   393 => x"ec050d76",
   394 => x"54805287",
   395 => x"0b881580",
   396 => x"f52d5653",
   397 => x"74722483",
   398 => x"38a05372",
   399 => x"5182f82d",
   400 => x"81128b15",
   401 => x"80f52d54",
   402 => x"52727225",
   403 => x"de380294",
   404 => x"050d0402",
   405 => x"f0050dac",
   406 => x"bc085481",
   407 => x"f72d800b",
   408 => x"acc00c73",
   409 => x"08802e81",
   410 => x"8038820b",
   411 => x"ac800cac",
   412 => x"c0088f06",
   413 => x"abfc0c73",
   414 => x"08527183",
   415 => x"2e963871",
   416 => x"83268938",
   417 => x"71812eaf",
   418 => x"388dd404",
   419 => x"71852e9f",
   420 => x"388dd404",
   421 => x"881480f5",
   422 => x"2d841508",
   423 => x"a8945354",
   424 => x"52859b2d",
   425 => x"71842913",
   426 => x"70085252",
   427 => x"8dd80473",
   428 => x"518ca32d",
   429 => x"8dd404ab",
   430 => x"bc088815",
   431 => x"082c7081",
   432 => x"06515271",
   433 => x"802e8738",
   434 => x"a898518d",
   435 => x"d104a89c",
   436 => x"51859b2d",
   437 => x"84140851",
   438 => x"859b2dac",
   439 => x"c0088105",
   440 => x"acc00c8c",
   441 => x"14548ce3",
   442 => x"04029005",
   443 => x"0d0471ac",
   444 => x"bc0c8cd3",
   445 => x"2dacc008",
   446 => x"ff05acc4",
   447 => x"0c0402e8",
   448 => x"050dacbc",
   449 => x"08acc808",
   450 => x"575580f6",
   451 => x"5189ad2d",
   452 => x"abec0881",
   453 => x"2a708106",
   454 => x"51527180",
   455 => x"2e9f388e",
   456 => x"a50487f6",
   457 => x"2d80f651",
   458 => x"89ad2dab",
   459 => x"ec08f338",
   460 => x"abe80881",
   461 => x"3270abe8",
   462 => x"0c51848a",
   463 => x"2d800bac",
   464 => x"b80c8c51",
   465 => x"89ad2dab",
   466 => x"ec08812a",
   467 => x"70810651",
   468 => x"5271802e",
   469 => x"bd38abc0",
   470 => x"08abd408",
   471 => x"abc00cab",
   472 => x"d40cabc4",
   473 => x"08abd808",
   474 => x"abc40cab",
   475 => x"d80cabc8",
   476 => x"08abdc08",
   477 => x"abc80cab",
   478 => x"dc0cabcc",
   479 => x"08abe008",
   480 => x"abcc0cab",
   481 => x"e00cabd0",
   482 => x"08abe408",
   483 => x"abd00cab",
   484 => x"e40cacb0",
   485 => x"08a00652",
   486 => x"80722594",
   487 => x"388bbb2d",
   488 => x"87f62dab",
   489 => x"e8088132",
   490 => x"70abe80c",
   491 => x"51848a2d",
   492 => x"abe80881",
   493 => x"ea38abd4",
   494 => x"085189ad",
   495 => x"2dabec08",
   496 => x"802e8938",
   497 => x"acb80881",
   498 => x"07acb80c",
   499 => x"abd80851",
   500 => x"89ad2dab",
   501 => x"ec08802e",
   502 => x"8938acb8",
   503 => x"088207ac",
   504 => x"b80cabdc",
   505 => x"085189ad",
   506 => x"2dabec08",
   507 => x"802e8938",
   508 => x"acb80884",
   509 => x"07acb80c",
   510 => x"abe00851",
   511 => x"89ad2dab",
   512 => x"ec08802e",
   513 => x"8938acb8",
   514 => x"088807ac",
   515 => x"b80cabe4",
   516 => x"085189ad",
   517 => x"2dabec08",
   518 => x"802e8938",
   519 => x"acb80890",
   520 => x"07acb80c",
   521 => x"abc00851",
   522 => x"89ad2dab",
   523 => x"ec08802e",
   524 => x"8a38acb8",
   525 => x"08828007",
   526 => x"acb80cab",
   527 => x"c4085189",
   528 => x"ad2dabec",
   529 => x"08802e8a",
   530 => x"38acb808",
   531 => x"848007ac",
   532 => x"b80cabc8",
   533 => x"085189ad",
   534 => x"2dabec08",
   535 => x"802e8a38",
   536 => x"acb80888",
   537 => x"8007acb8",
   538 => x"0cabcc08",
   539 => x"5189ad2d",
   540 => x"abec0880",
   541 => x"2e8a38ac",
   542 => x"b8089080",
   543 => x"07acb80c",
   544 => x"abd00851",
   545 => x"89ad2dab",
   546 => x"ec08802e",
   547 => x"8a38acb8",
   548 => x"08a08007",
   549 => x"acb80cac",
   550 => x"b808ed0c",
   551 => x"97fc04ab",
   552 => x"e4085189",
   553 => x"ad2dabec",
   554 => x"08802e89",
   555 => x"38acb808",
   556 => x"9007acb8",
   557 => x"0cacb808",
   558 => x"ed0c81f5",
   559 => x"5189ad2d",
   560 => x"abec0881",
   561 => x"2a708106",
   562 => x"515271a0",
   563 => x"38abd408",
   564 => x"5189ad2d",
   565 => x"abec0881",
   566 => x"2a708106",
   567 => x"5152718c",
   568 => x"38acb008",
   569 => x"90065280",
   570 => x"7225bd38",
   571 => x"acb00890",
   572 => x"06528072",
   573 => x"2584388b",
   574 => x"bb2dacc4",
   575 => x"08527180",
   576 => x"2e8938ff",
   577 => x"12acc40c",
   578 => x"92a804ac",
   579 => x"c00810ac",
   580 => x"c0080570",
   581 => x"84291651",
   582 => x"52881208",
   583 => x"802e8938",
   584 => x"ff518812",
   585 => x"0852712d",
   586 => x"81f25189",
   587 => x"ad2dabec",
   588 => x"08812a70",
   589 => x"81065152",
   590 => x"71a038ab",
   591 => x"d8085189",
   592 => x"ad2dabec",
   593 => x"08812a70",
   594 => x"81065152",
   595 => x"718c38ac",
   596 => x"b0088806",
   597 => x"52807225",
   598 => x"bf38acb0",
   599 => x"08880652",
   600 => x"80722584",
   601 => x"388bbb2d",
   602 => x"acc008ff",
   603 => x"11acc408",
   604 => x"56535373",
   605 => x"72258938",
   606 => x"8114acc4",
   607 => x"0c939804",
   608 => x"72101370",
   609 => x"84291651",
   610 => x"52881208",
   611 => x"802e8938",
   612 => x"fe518812",
   613 => x"0852712d",
   614 => x"81fd5189",
   615 => x"ad2dabec",
   616 => x"08812a70",
   617 => x"81065152",
   618 => x"719738ab",
   619 => x"dc085189",
   620 => x"ad2dabec",
   621 => x"08812a70",
   622 => x"81065152",
   623 => x"71802ead",
   624 => x"38acc408",
   625 => x"802e8938",
   626 => x"800bacc4",
   627 => x"0c93ed04",
   628 => x"acc00810",
   629 => x"acc00805",
   630 => x"70842916",
   631 => x"51528812",
   632 => x"08802e89",
   633 => x"38fd5188",
   634 => x"12085271",
   635 => x"2d81fa51",
   636 => x"89ad2dab",
   637 => x"ec08812a",
   638 => x"70810651",
   639 => x"52719738",
   640 => x"abe00851",
   641 => x"89ad2dab",
   642 => x"ec08812a",
   643 => x"70810651",
   644 => x"5271802e",
   645 => x"ae38acc0",
   646 => x"08ff1154",
   647 => x"52acc408",
   648 => x"73258838",
   649 => x"72acc40c",
   650 => x"94c30471",
   651 => x"10127084",
   652 => x"29165152",
   653 => x"88120880",
   654 => x"2e8938fc",
   655 => x"51881208",
   656 => x"52712dac",
   657 => x"c4087053",
   658 => x"5473802e",
   659 => x"8a388c15",
   660 => x"ff155555",
   661 => x"94c90482",
   662 => x"0bac800c",
   663 => x"718f06ab",
   664 => x"fc0c81eb",
   665 => x"5189ad2d",
   666 => x"abec0881",
   667 => x"2a708106",
   668 => x"51527180",
   669 => x"2ead3874",
   670 => x"08852e09",
   671 => x"8106a438",
   672 => x"881580f5",
   673 => x"2dff0552",
   674 => x"71881681",
   675 => x"b72d7198",
   676 => x"2b527180",
   677 => x"25883880",
   678 => x"0b881681",
   679 => x"b72d7451",
   680 => x"8ca32d81",
   681 => x"f45189ad",
   682 => x"2dabec08",
   683 => x"812a7081",
   684 => x"06515271",
   685 => x"802eb338",
   686 => x"7408852e",
   687 => x"098106aa",
   688 => x"38881580",
   689 => x"f52d8105",
   690 => x"52718816",
   691 => x"81b72d71",
   692 => x"81ff068b",
   693 => x"1680f52d",
   694 => x"54527272",
   695 => x"27873872",
   696 => x"881681b7",
   697 => x"2d74518c",
   698 => x"a32d80da",
   699 => x"5189ad2d",
   700 => x"abec0881",
   701 => x"2a708106",
   702 => x"5152718d",
   703 => x"38acb008",
   704 => x"81065280",
   705 => x"722581b4",
   706 => x"38acbc08",
   707 => x"acb00881",
   708 => x"06535380",
   709 => x"72258438",
   710 => x"8bbb2dac",
   711 => x"c4085473",
   712 => x"802e8a38",
   713 => x"8c13ff15",
   714 => x"5553969f",
   715 => x"04720852",
   716 => x"71822ea6",
   717 => x"38718226",
   718 => x"89387181",
   719 => x"2ea93897",
   720 => x"bc047183",
   721 => x"2eb13871",
   722 => x"842e0981",
   723 => x"0680ed38",
   724 => x"88130851",
   725 => x"8dee2d97",
   726 => x"bc04acc4",
   727 => x"08518813",
   728 => x"0852712d",
   729 => x"97bc0481",
   730 => x"0b881408",
   731 => x"2babbc08",
   732 => x"32abbc0c",
   733 => x"97920488",
   734 => x"1380f52d",
   735 => x"81058b14",
   736 => x"80f52d53",
   737 => x"54717424",
   738 => x"83388054",
   739 => x"73881481",
   740 => x"b72d8cd3",
   741 => x"2d97bc04",
   742 => x"7508802e",
   743 => x"a2387508",
   744 => x"5189ad2d",
   745 => x"abec0881",
   746 => x"06527180",
   747 => x"2e8b38ac",
   748 => x"c4085184",
   749 => x"16085271",
   750 => x"2d881656",
   751 => x"75da3880",
   752 => x"54800bac",
   753 => x"800c738f",
   754 => x"06abfc0c",
   755 => x"a05273ac",
   756 => x"c4082e09",
   757 => x"81069838",
   758 => x"acc008ff",
   759 => x"05743270",
   760 => x"09810570",
   761 => x"72079f2a",
   762 => x"91713151",
   763 => x"51535371",
   764 => x"5182f82d",
   765 => x"8114548e",
   766 => x"7425c638",
   767 => x"abe808ab",
   768 => x"ec0c0298",
   769 => x"050d0402",
   770 => x"f4050dd4",
   771 => x"5281ff72",
   772 => x"0c710853",
   773 => x"81ff720c",
   774 => x"72882b83",
   775 => x"fe800672",
   776 => x"087081ff",
   777 => x"06515253",
   778 => x"81ff720c",
   779 => x"72710788",
   780 => x"2b720870",
   781 => x"81ff0651",
   782 => x"525381ff",
   783 => x"720c7271",
   784 => x"07882b72",
   785 => x"087081ff",
   786 => x"067207ab",
   787 => x"ec0c5253",
   788 => x"028c050d",
   789 => x"0402f405",
   790 => x"0d747671",
   791 => x"81ff06d4",
   792 => x"0c5353ac",
   793 => x"cc088538",
   794 => x"71892b52",
   795 => x"71982ad4",
   796 => x"0c71902a",
   797 => x"7081ff06",
   798 => x"d40c5171",
   799 => x"882a7081",
   800 => x"ff06d40c",
   801 => x"517181ff",
   802 => x"06d40c72",
   803 => x"902a7081",
   804 => x"ff06d40c",
   805 => x"51d40870",
   806 => x"81ff0651",
   807 => x"5182b8bf",
   808 => x"527081ff",
   809 => x"2e098106",
   810 => x"943881ff",
   811 => x"0bd40cd4",
   812 => x"087081ff",
   813 => x"06ff1454",
   814 => x"515171e5",
   815 => x"3870abec",
   816 => x"0c028c05",
   817 => x"0d0402fc",
   818 => x"050d81c7",
   819 => x"5181ff0b",
   820 => x"d40cff11",
   821 => x"51708025",
   822 => x"f4380284",
   823 => x"050d0402",
   824 => x"f4050d81",
   825 => x"ff0bd40c",
   826 => x"93538052",
   827 => x"87fc80c1",
   828 => x"5198d52d",
   829 => x"abec088b",
   830 => x"3881ff0b",
   831 => x"d40c8153",
   832 => x"9a8c0499",
   833 => x"c62dff13",
   834 => x"5372df38",
   835 => x"72abec0c",
   836 => x"028c050d",
   837 => x"0402ec05",
   838 => x"0d810bac",
   839 => x"cc0c8454",
   840 => x"d008708f",
   841 => x"2a708106",
   842 => x"51515372",
   843 => x"f33872d0",
   844 => x"0c99c62d",
   845 => x"a8a05185",
   846 => x"9b2dd008",
   847 => x"708f2a70",
   848 => x"81065151",
   849 => x"5372f338",
   850 => x"810bd00c",
   851 => x"b1538052",
   852 => x"84d480c0",
   853 => x"5198d52d",
   854 => x"abec0881",
   855 => x"2e933872",
   856 => x"822ebd38",
   857 => x"ff135372",
   858 => x"e538ff14",
   859 => x"5473ffb0",
   860 => x"3899c62d",
   861 => x"83aa5284",
   862 => x"9c80c851",
   863 => x"98d52dab",
   864 => x"ec08812e",
   865 => x"09810692",
   866 => x"3898872d",
   867 => x"abec0883",
   868 => x"ffff0653",
   869 => x"7283aa2e",
   870 => x"9d3899df",
   871 => x"2d9bb104",
   872 => x"a8ac5185",
   873 => x"9b2d8053",
   874 => x"9cff04a8",
   875 => x"c451859b",
   876 => x"2d80549c",
   877 => x"d10481ff",
   878 => x"0bd40cb1",
   879 => x"5499c62d",
   880 => x"8fcf5380",
   881 => x"5287fc80",
   882 => x"f75198d5",
   883 => x"2dabec08",
   884 => x"55abec08",
   885 => x"812e0981",
   886 => x"069b3881",
   887 => x"ff0bd40c",
   888 => x"820a5284",
   889 => x"9c80e951",
   890 => x"98d52dab",
   891 => x"ec08802e",
   892 => x"8d3899c6",
   893 => x"2dff1353",
   894 => x"72c9389c",
   895 => x"c40481ff",
   896 => x"0bd40cab",
   897 => x"ec085287",
   898 => x"fc80fa51",
   899 => x"98d52dab",
   900 => x"ec08b138",
   901 => x"81ff0bd4",
   902 => x"0cd40853",
   903 => x"81ff0bd4",
   904 => x"0c81ff0b",
   905 => x"d40c81ff",
   906 => x"0bd40c81",
   907 => x"ff0bd40c",
   908 => x"72862a70",
   909 => x"81067656",
   910 => x"51537295",
   911 => x"38abec08",
   912 => x"549cd104",
   913 => x"73822efe",
   914 => x"e238ff14",
   915 => x"5473feed",
   916 => x"3873accc",
   917 => x"0c738b38",
   918 => x"815287fc",
   919 => x"80d05198",
   920 => x"d52d81ff",
   921 => x"0bd40cd0",
   922 => x"08708f2a",
   923 => x"70810651",
   924 => x"515372f3",
   925 => x"3872d00c",
   926 => x"81ff0bd4",
   927 => x"0c815372",
   928 => x"abec0c02",
   929 => x"94050d04",
   930 => x"02e8050d",
   931 => x"78558056",
   932 => x"81ff0bd4",
   933 => x"0cd00870",
   934 => x"8f2a7081",
   935 => x"06515153",
   936 => x"72f33882",
   937 => x"810bd00c",
   938 => x"81ff0bd4",
   939 => x"0c775287",
   940 => x"fc80d151",
   941 => x"98d52d80",
   942 => x"dbc6df54",
   943 => x"abec0880",
   944 => x"2e8a38a8",
   945 => x"e451859b",
   946 => x"2d9e9f04",
   947 => x"81ff0bd4",
   948 => x"0cd40870",
   949 => x"81ff0651",
   950 => x"537281fe",
   951 => x"2e098106",
   952 => x"9d3880ff",
   953 => x"5398872d",
   954 => x"abec0875",
   955 => x"70840557",
   956 => x"0cff1353",
   957 => x"728025ed",
   958 => x"3881569e",
   959 => x"8404ff14",
   960 => x"5473c938",
   961 => x"81ff0bd4",
   962 => x"0c81ff0b",
   963 => x"d40cd008",
   964 => x"708f2a70",
   965 => x"81065151",
   966 => x"5372f338",
   967 => x"72d00c75",
   968 => x"abec0c02",
   969 => x"98050d04",
   970 => x"02e8050d",
   971 => x"77797b58",
   972 => x"55558053",
   973 => x"727625a3",
   974 => x"38747081",
   975 => x"055680f5",
   976 => x"2d747081",
   977 => x"055680f5",
   978 => x"2d525271",
   979 => x"712e8638",
   980 => x"81519edd",
   981 => x"04811353",
   982 => x"9eb40480",
   983 => x"5170abec",
   984 => x"0c029805",
   985 => x"0d0402ec",
   986 => x"050d7655",
   987 => x"74802ebb",
   988 => x"389a1580",
   989 => x"e02d51a5",
   990 => x"ea2dabec",
   991 => x"08abec08",
   992 => x"b0fc0cab",
   993 => x"ec085454",
   994 => x"b0d80880",
   995 => x"2e993894",
   996 => x"1580e02d",
   997 => x"51a5ea2d",
   998 => x"abec0890",
   999 => x"2b83fff0",
  1000 => x"0a067075",
  1001 => x"07515372",
  1002 => x"b0fc0cb0",
  1003 => x"fc085372",
  1004 => x"802e9938",
  1005 => x"b0d008fe",
  1006 => x"147129b0",
  1007 => x"e40805b1",
  1008 => x"800c7084",
  1009 => x"2bb0dc0c",
  1010 => x"549ff204",
  1011 => x"b0e808b0",
  1012 => x"fc0cb0ec",
  1013 => x"08b1800c",
  1014 => x"b0d80880",
  1015 => x"2e8a38b0",
  1016 => x"d008842b",
  1017 => x"539fee04",
  1018 => x"b0f00884",
  1019 => x"2b5372b0",
  1020 => x"dc0c0294",
  1021 => x"050d0402",
  1022 => x"d8050d80",
  1023 => x"0bb0d80c",
  1024 => x"84549a95",
  1025 => x"2dabec08",
  1026 => x"802e9538",
  1027 => x"acd05280",
  1028 => x"519d882d",
  1029 => x"abec0880",
  1030 => x"2e8638fe",
  1031 => x"54a0a804",
  1032 => x"ff145473",
  1033 => x"8024db38",
  1034 => x"738c38a8",
  1035 => x"f451859b",
  1036 => x"2d7355a5",
  1037 => x"b1048056",
  1038 => x"810bb184",
  1039 => x"0c8853a9",
  1040 => x"8852ad86",
  1041 => x"519ea82d",
  1042 => x"abec0876",
  1043 => x"2e098106",
  1044 => x"8738abec",
  1045 => x"08b1840c",
  1046 => x"8853a994",
  1047 => x"52ada251",
  1048 => x"9ea82dab",
  1049 => x"ec088738",
  1050 => x"abec08b1",
  1051 => x"840cb184",
  1052 => x"08802e80",
  1053 => x"f638b096",
  1054 => x"0b80f52d",
  1055 => x"b0970b80",
  1056 => x"f52d7198",
  1057 => x"2b71902b",
  1058 => x"07b0980b",
  1059 => x"80f52d70",
  1060 => x"882b7207",
  1061 => x"b0990b80",
  1062 => x"f52d7107",
  1063 => x"b0ce0b80",
  1064 => x"f52db0cf",
  1065 => x"0b80f52d",
  1066 => x"71882b07",
  1067 => x"535f5452",
  1068 => x"5a565755",
  1069 => x"7381abaa",
  1070 => x"2e098106",
  1071 => x"8d387551",
  1072 => x"a5ba2dab",
  1073 => x"ec0856a1",
  1074 => x"d7047382",
  1075 => x"d4d52e87",
  1076 => x"38a9a051",
  1077 => x"a29804ac",
  1078 => x"d0527551",
  1079 => x"9d882dab",
  1080 => x"ec0855ab",
  1081 => x"ec08802e",
  1082 => x"83c73888",
  1083 => x"53a99452",
  1084 => x"ada2519e",
  1085 => x"a82dabec",
  1086 => x"08893881",
  1087 => x"0bb0d80c",
  1088 => x"a29e0488",
  1089 => x"53a98852",
  1090 => x"ad86519e",
  1091 => x"a82dabec",
  1092 => x"08802e8a",
  1093 => x"38a9b451",
  1094 => x"859b2da2",
  1095 => x"f804b0ce",
  1096 => x"0b80f52d",
  1097 => x"547380d5",
  1098 => x"2e098106",
  1099 => x"80ca38b0",
  1100 => x"cf0b80f5",
  1101 => x"2d547381",
  1102 => x"aa2e0981",
  1103 => x"06ba3880",
  1104 => x"0bacd00b",
  1105 => x"80f52d56",
  1106 => x"547481e9",
  1107 => x"2e833881",
  1108 => x"547481eb",
  1109 => x"2e8c3880",
  1110 => x"5573752e",
  1111 => x"09810682",
  1112 => x"d038acdb",
  1113 => x"0b80f52d",
  1114 => x"55748d38",
  1115 => x"acdc0b80",
  1116 => x"f52d5473",
  1117 => x"822e8638",
  1118 => x"8055a5b1",
  1119 => x"04acdd0b",
  1120 => x"80f52d70",
  1121 => x"b0d00cff",
  1122 => x"05b0d40c",
  1123 => x"acde0b80",
  1124 => x"f52dacdf",
  1125 => x"0b80f52d",
  1126 => x"58760577",
  1127 => x"82802905",
  1128 => x"70b0e00c",
  1129 => x"ace00b80",
  1130 => x"f52d70b0",
  1131 => x"f40cb0d8",
  1132 => x"08595758",
  1133 => x"76802e81",
  1134 => x"a3388853",
  1135 => x"a99452ad",
  1136 => x"a2519ea8",
  1137 => x"2dabec08",
  1138 => x"81e738b0",
  1139 => x"d0087084",
  1140 => x"2bb0dc0c",
  1141 => x"70b0f00c",
  1142 => x"acf50b80",
  1143 => x"f52dacf4",
  1144 => x"0b80f52d",
  1145 => x"71828029",
  1146 => x"05acf60b",
  1147 => x"80f52d70",
  1148 => x"84808029",
  1149 => x"12acf70b",
  1150 => x"80f52d70",
  1151 => x"81800a29",
  1152 => x"1270b0f8",
  1153 => x"0cb0f408",
  1154 => x"7129b0e0",
  1155 => x"080570b0",
  1156 => x"e40cacfd",
  1157 => x"0b80f52d",
  1158 => x"acfc0b80",
  1159 => x"f52d7182",
  1160 => x"802905ac",
  1161 => x"fe0b80f5",
  1162 => x"2d708480",
  1163 => x"802912ac",
  1164 => x"ff0b80f5",
  1165 => x"2d70982b",
  1166 => x"81f00a06",
  1167 => x"720570b0",
  1168 => x"e80cfe11",
  1169 => x"7e297705",
  1170 => x"b0ec0c52",
  1171 => x"59524354",
  1172 => x"5e515259",
  1173 => x"525d5759",
  1174 => x"57a5aa04",
  1175 => x"ace20b80",
  1176 => x"f52dace1",
  1177 => x"0b80f52d",
  1178 => x"71828029",
  1179 => x"0570b0dc",
  1180 => x"0c70a029",
  1181 => x"83ff0570",
  1182 => x"892a70b0",
  1183 => x"f00cace7",
  1184 => x"0b80f52d",
  1185 => x"ace60b80",
  1186 => x"f52d7182",
  1187 => x"80290570",
  1188 => x"b0f80c7b",
  1189 => x"71291e70",
  1190 => x"b0ec0c7d",
  1191 => x"b0e80c73",
  1192 => x"05b0e40c",
  1193 => x"555e5151",
  1194 => x"55558051",
  1195 => x"9ee62d81",
  1196 => x"5574abec",
  1197 => x"0c02a805",
  1198 => x"0d0402f4",
  1199 => x"050d7470",
  1200 => x"882a83fe",
  1201 => x"80067072",
  1202 => x"982a0772",
  1203 => x"882b87fc",
  1204 => x"80800673",
  1205 => x"982b81f0",
  1206 => x"0a067173",
  1207 => x"0707abec",
  1208 => x"0c565153",
  1209 => x"51028c05",
  1210 => x"0d0402f8",
  1211 => x"050d028e",
  1212 => x"0580f52d",
  1213 => x"74882b07",
  1214 => x"7083ffff",
  1215 => x"06abec0c",
  1216 => x"51028805",
  1217 => x"0d040000",
  1218 => x"00ffffff",
  1219 => x"ff00ffff",
  1220 => x"ffff00ff",
  1221 => x"ffffff00",
  1222 => x"52657365",
  1223 => x"74000000",
  1224 => x"4d616e75",
  1225 => x"616c2053",
  1226 => x"65727665",
  1227 => x"00000000",
  1228 => x"42616c6c",
  1229 => x"20416e67",
  1230 => x"6c650000",
  1231 => x"42616c6c",
  1232 => x"20537065",
  1233 => x"65640000",
  1234 => x"50616464",
  1235 => x"6c652053",
  1236 => x"697a6500",
  1237 => x"536f756e",
  1238 => x"64000000",
  1239 => x"466f7572",
  1240 => x"20706c61",
  1241 => x"79657273",
  1242 => x"00000000",
  1243 => x"446f7562",
  1244 => x"6c65204f",
  1245 => x"53442077",
  1246 => x"696e646f",
  1247 => x"77000000",
  1248 => x"45786974",
  1249 => x"00000000",
  1250 => x"4d6f6e6f",
  1251 => x"00000000",
  1252 => x"47726579",
  1253 => x"7363616c",
  1254 => x"65000000",
  1255 => x"52474231",
  1256 => x"00000000",
  1257 => x"52474232",
  1258 => x"00000000",
  1259 => x"4669656c",
  1260 => x"64000000",
  1261 => x"49636500",
  1262 => x"43687269",
  1263 => x"73746d61",
  1264 => x"73000000",
  1265 => x"4d61726b",
  1266 => x"736d616e",
  1267 => x"00000000",
  1268 => x"4c617320",
  1269 => x"56656761",
  1270 => x"73000000",
  1271 => x"41592d33",
  1272 => x"2d383531",
  1273 => x"3520636f",
  1274 => x"6c6f7273",
  1275 => x"00000000",
  1276 => x"54525120",
  1277 => x"436f6c6f",
  1278 => x"72730000",
  1279 => x"496e6974",
  1280 => x"69616c69",
  1281 => x"7a696e67",
  1282 => x"20534420",
  1283 => x"63617264",
  1284 => x"0a000000",
  1285 => x"16200000",
  1286 => x"14200000",
  1287 => x"15200000",
  1288 => x"53442069",
  1289 => x"6e69742e",
  1290 => x"2e2e0a00",
  1291 => x"53442063",
  1292 => x"61726420",
  1293 => x"72657365",
  1294 => x"74206661",
  1295 => x"696c6564",
  1296 => x"210a0000",
  1297 => x"53444843",
  1298 => x"20657272",
  1299 => x"6f72210a",
  1300 => x"00000000",
  1301 => x"57726974",
  1302 => x"65206661",
  1303 => x"696c6564",
  1304 => x"0a000000",
  1305 => x"52656164",
  1306 => x"20666169",
  1307 => x"6c65640a",
  1308 => x"00000000",
  1309 => x"43617264",
  1310 => x"20696e69",
  1311 => x"74206661",
  1312 => x"696c6564",
  1313 => x"0a000000",
  1314 => x"46415431",
  1315 => x"36202020",
  1316 => x"00000000",
  1317 => x"46415433",
  1318 => x"32202020",
  1319 => x"00000000",
  1320 => x"4e6f2070",
  1321 => x"61727469",
  1322 => x"74696f6e",
  1323 => x"20736967",
  1324 => x"0a000000",
  1325 => x"42616420",
  1326 => x"70617274",
  1327 => x"0a000000",
  1328 => x"00000002",
  1329 => x"00000002",
  1330 => x"00001318",
  1331 => x"000002d4",
  1332 => x"00000001",
  1333 => x"00001320",
  1334 => x"00000000",
  1335 => x"00000001",
  1336 => x"00001330",
  1337 => x"00000001",
  1338 => x"00000001",
  1339 => x"0000133c",
  1340 => x"00000002",
  1341 => x"00000001",
  1342 => x"00001348",
  1343 => x"00000003",
  1344 => x"00000001",
  1345 => x"00001354",
  1346 => x"00000004",
  1347 => x"00000001",
  1348 => x"0000135c",
  1349 => x"00000006",
  1350 => x"00000001",
  1351 => x"0000136c",
  1352 => x"00000005",
  1353 => x"00000003",
  1354 => x"00001548",
  1355 => x"0000000b",
  1356 => x"00000002",
  1357 => x"00001380",
  1358 => x"000005e5",
  1359 => x"00000000",
  1360 => x"00000000",
  1361 => x"00000000",
  1362 => x"00001388",
  1363 => x"00001390",
  1364 => x"0000139c",
  1365 => x"000013a4",
  1366 => x"000013ac",
  1367 => x"000013b4",
  1368 => x"000013b8",
  1369 => x"000013c4",
  1370 => x"000013d0",
  1371 => x"000013dc",
  1372 => x"000013f0",
  1373 => x"00000000",
  1374 => x"00000000",
  1375 => x"00000000",
  1376 => x"00000000",
  1377 => x"00000000",
  1378 => x"00000000",
  1379 => x"00000000",
  1380 => x"00000000",
  1381 => x"00000000",
  1382 => x"00000000",
  1383 => x"00000000",
  1384 => x"00000000",
  1385 => x"00000000",
  1386 => x"00000000",
  1387 => x"00000000",
  1388 => x"00000000",
  1389 => x"00000000",
  1390 => x"00000000",
  1391 => x"00000006",
  1392 => x"00000043",
  1393 => x"00000042",
  1394 => x"0000003b",
  1395 => x"0000004b",
  1396 => x"0000007e",
  1397 => x"00000003",
  1398 => x"0000000b",
  1399 => x"00000083",
  1400 => x"00000023",
  1401 => x"0000007e",
  1402 => x"00000000",
	others => x"00000000"
);

begin

process (clk)
begin
	if (clk'event and clk = '1') then
		if (from_zpu.memAWriteEnable = '1') and (from_zpu.memBWriteEnable = '1') and (from_zpu.memAAddr=from_zpu.memBAddr) and (from_zpu.memAWrite/=from_zpu.memBWrite) then
			report "write collision" severity failure;
		end if;
	
		if (from_zpu.memAWriteEnable = '1') then
			ram(to_integer(unsigned(from_zpu.memAAddr(maxAddrBitBRAM downto 2)))) := from_zpu.memAWrite;
			to_zpu.memARead <= from_zpu.memAWrite;
		else
			to_zpu.memARead <= ram(to_integer(unsigned(from_zpu.memAAddr(maxAddrBitBRAM downto 2))));
		end if;
	end if;
end process;

process (clk)
begin
	if (clk'event and clk = '1') then
		if (from_zpu.memBWriteEnable = '1') then
			ram(to_integer(unsigned(from_zpu.memBAddr(maxAddrBitBRAM downto 2)))) := from_zpu.memBWrite;
			to_zpu.memBRead <= from_zpu.memBWrite;
		else
			to_zpu.memBRead <= ram(to_integer(unsigned(from_zpu.memBAddr(maxAddrBitBRAM downto 2))));
		end if;
	end if;
end process;


end arch;

