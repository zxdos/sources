00
ff
00
e0
60
00
61
38
68
00
69
00
6a
00
6b
00
6c
7f
6d
32
a3
6c
d0
12
70
08
40
80
12
20
12
16
23
30
23
58
60
0e
e0
a1
12
34
60
0f
e0
a1
12
38
12
24
12
32
66
01
12
3a
66
00
86
60
60
01
f0
18
60
01
f0
15
f0
07
30
00
12
44
60
01
e0
a1
23
18
60
04
e0
a1
23
24
60
02
e0
a1
22
b8
46
01
12
d8
60
0c
e0
a1
23
00
60
0d
e0
a1
23
0c
60
03
e0
a1
22
74
12
e6
a3
60
60
00
d0
d6
84
f0
60
05
f0
18
60
00
d0
d6
44
01
12
8a
00
ee
23
30
79
01
23
30
49
63
12
32
00
ee
a3
60
60
00
d0
d6
84
f0
60
05
f0
18
60
00
d0
d6
44
01
12
ac
12
e6
23
30
79
01
23
30
49
63
12
32
12
e6
60
7f
d0
b6
60
05
f0
18
84
f0
60
7f
d0
b6
44
01
12
cc
00
ee
23
30
78
01
23
30
48
63
12
32
00
ee
c0
03
40
00
12
96
40
01
12
e8
40
02
12
f4
12
3c
4d
00
12
e6
23
58
7d
fe
23
58
12
e6
4d
32
12
e6
23
58
7d
02
23
58
12
e6
4d
00
00
ee
23
58
7d
fe
23
58
00
ee
4d
32
00
ee
23
58
7d
02
23
58
00
ee
4b
00
00
ee
23
58
7b
fe
23
58
00
ee
4b
32
00
ee
23
58
7b
02
23
58
00
ee
a3
66
63
00
64
3b
f8
33
f2
65
f1
29
d3
45
73
05
f2
29
d3
45
63
77
a3
66
f9
33
f2
65
f1
29
d3
45
f2
29
73
05
d3
45
00
ee
a3
60
da
b6
dc
d6
00
ee
80
80
80
80
80
80
00
00
00
00
00
00
ff
ff
