12
0e
5b
20
41
6e
74
20
76
31
2e
30
20
5d
00
ff
60
fe
61
00
aa
10
f1
55
22
4c
23
5c
65
00
6a
01
6b
00
6d
00
6e
00
23
68
3f
00
13
c6
45
fd
12
d0
47
cc
22
7a
41
fb
14
d0
41
fc
15
68
41
fa
15
e0
41
f9
16
2c
60
02
37
cc
24
c6
12
26
6e
00
a7
f2
fe
1e
60
2e
f0
55
70
09
61
7c
aa
e8
d1
04
60
01
24
c0
60
02
24
c6
3e
1f
00
fc
7e
01
3e
20
12
4e
60
04
61
04
aa
f8
d0
10
00
ee
4b
00
22
e6
7b
ff
aa
12
f1
65
a7
f2
fe
1e
f0
55
7e
01
62
1f
8e
22
41
fe
12
a4
41
ff
12
ae
70
09
62
7c
aa
e8
fd
1e
d2
04
00
ee
70
07
61
7c
ab
38
d1
04
00
ee
61
00
4b
02
61
08
4b
01
61
10
4b
00
61
18
ab
18
f1
1e
61
7c
70
01
d1
08
70
08
aa
e8
fd
1e
d1
04
00
ee
47
cc
73
fc
ad
5c
d3
40
33
00
73
fc
33
00
d3
40
43
00
65
00
12
30
aa
10
f1
65
70
02
40
fe
23
1a
f0
55
a8
12
41
01
a9
10
f0
1e
f1
65
aa
12
f1
55
62
f0
82
17
4f
00
13
16
41
fe
13
24
41
ff
13
28
41
fd
13
2c
13
58
8b
10
00
ee
61
01
60
00
aa
10
f1
55
00
ee
6b
0c
00
ee
6b
04
00
ee
6b
01
65
fd
84
00
74
f9
60
70
ab
dc
d0
40
60
04
24
c0
63
60
ad
5c
d3
40
60
02
24
c0
60
02
24
c6
60
01
24
c0
60
70
ab
dc
d0
40
00
ee
6b
01
00
ee
66
00
68
2e
6c
00
aa
68
d6
80
00
ee
67
00
24
2e
23
de
82
c0
60
0c
e0
a1
24
66
60
03
e0
a1
24
86
80
60
37
cc
86
74
81
80
88
94
aa
68
f2
1e
d0
10
47
cc
00
fc
aa
68
fc
1e
d6
80
00
ee
67
00
24
2e
23
de
82
c0
60
0c
e0
a1
24
66
47
cc
67
04
60
03
e0
a1
24
86
80
60
86
74
81
80
88
94
aa
68
f2
1e
d0
10
aa
68
fc
1e
d6
80
00
ee
61
00
d6
80
60
02
24
c0
60
02
24
c6
71
01
31
07
13
c8
60
1e
24
c6
00
fd
60
0a
e0
9e
14
0c
4a
00
00
ee
4a
01
23
fe
6a
02
69
fc
aa
0e
f0
65
58
00
00
ee
6a
00
69
fe
00
ee
60
02
24
c0
80
80
70
ec
aa
0e
f0
55
00
ee
4a
02
14
28
80
60
24
52
98
00
14
24
80
60
70
0c
24
52
98
00
14
24
00
ee
6a
01
00
ee
6a
00
69
fe
00
ee
4a
02
00
ee
60
04
49
fe
60
02
89
00
80
60
24
52
98
00
69
00
80
60
70
0c
24
52
98
00
69
00
49
04
6a
00
00
ee
80
56
80
56
80
e4
61
1f
80
12
a7
f2
f0
1e
f0
65
81
00
00
ee
60
00
4c
00
60
20
8c
00
80
60
70
10
24
52
80
85
4f
00
00
ee
67
04
46
38
67
cc
91
80
14
b2
00
ee
60
40
4c
40
60
60
8c
00
46
00
00
ee
80
60
70
fc
24
52
80
85
4f
00
00
ee
67
fc
91
80
14
a6
00
ee
80
60
24
52
80
87
4f
00
69
fc
00
ee
80
60
70
0c
24
52
80
87
4f
00
69
fc
00
ee
f0
18
80
5e
14
c6
f0
15
f0
07
30
00
14
c8
00
ee
24
e2
24
f6
23
98
3f
00
13
c6
25
10
46
70
15
3c
14
d4
60
01
24
c0
aa
68
fc
1e
d6
80
76
fc
d6
80
36
00
14
e2
00
ee
63
09
64
25
65
04
60
18
ab
3c
d0
30
70
14
d0
40
70
14
d0
30
70
14
d0
40
00
ee
43
09
65
04
43
25
65
fc
ab
3c
60
18
81
30
83
54
d0
10
d0
30
60
40
d0
10
d0
30
60
2c
81
40
84
55
d0
10
d0
40
60
54
d0
10
d0
40
00
ee
7d
04
00
fc
a7
f2
fe
1e
60
2a
f0
55
70
09
61
7c
aa
e8
fd
1e
d1
04
60
01
24
c0
60
02
24
c6
7e
01
4e
20
6e
00
76
fc
36
00
15
3e
12
26
24
e2
25
7a
25
8c
23
98
3f
00
13
c6
46
70
15
3c
15
6c
60
70
61
0f
62
fe
63
00
aa
14
f3
55
ab
5c
d0
10
00
ee
aa
14
f3
65
84
20
42
02
64
fe
42
fe
64
02
41
11
25
cc
41
21
25
d4
82
40
84
30
73
20
43
80
63
00
ab
5c
f4
1e
84
10
81
24
85
00
70
fc
d5
40
ab
5c
f3
1e
35
00
d0
10
aa
14
f3
55
35
00
00
ee
15
7a
64
04
42
fc
64
fe
00
ee
64
fc
42
04
64
02
44
02
f4
18
00
ee
25
f0
25
fc
23
98
3f
00
13
c6
36
70
15
e2
15
3c
63
70
64
0f
65
00
ad
7c
d3
40
00
ee
80
30
70
0c
24
52
71
f9
54
10
26
22
80
30
73
fc
ad
7c
f5
1e
75
20
d0
10
ad
7c
f5
1e
30
00
d3
40
30
00
00
ee
15
f0
81
40
74
04
60
02
f0
18
00
ee
24
e2
26
5c
6e
00
26
68
27
48
3f
00
13
c6
46
70
17
d6
26
46
60
03
24
c6
16
34
4d
00
16
d0
4d
02
16
f6
4d
04
16
a8
4d
06
16
80
4d
08
17
2e
17
40
63
68
64
27
65
00
ab
dc
d3
40
00
ee
6b
00
65
00
aa
54
fe
1e
f0
65
8d
00
7e
01
4e
14
6e
00
4d
08
17
1c
00
ee
64
27
82
50
75
20
45
40
65
00
80
30
73
04
ac
dc
f2
1e
40
48
ab
dc
d0
40
ac
dc
f5
1e
43
68
ab
dc
d3
40
33
68
00
ee
16
68
64
27
82
50
75
20
45
40
65
00
80
30
73
fc
ad
1c
f2
1e
40
68
ab
dc
d0
40
ad
1c
f5
1e
43
48
ab
dc
d3
40
33
48
00
ee
16
68
aa
18
fb
1e
f2
65
ab
dc
f5
1e
d3
40
ab
dc
f2
1e
d0
10
83
00
84
10
85
20
60
01
45
20
24
c0
7b
03
3b
1e
00
ee
16
68
aa
36
fb
1e
f2
65
ab
dc
f5
1e
d3
40
ab
dc
f2
1e
d0
10
83
00
84
10
85
20
60
01
45
20
24
c0
7b
03
3b
1e
00
ee
16
68
85
30
75
f0
ad
5c
d5
40
60
01
24
c0
60
01
24
c0
00
ee
80
50
75
fc
ad
5c
d0
40
30
00
d5
40
30
00
00
ee
16
68
75
01
35
06
00
ee
16
68
67
00
27
a4
27
72
82
c0
60
0c
e0
a1
27
ba
60
03
e0
a1
27
c6
80
60
86
74
81
80
88
94
aa
68
f2
1e
d0
10
aa
68
fc
1e
d6
80
00
ee
60
0a
e0
9e
17
90
4a
00
00
ee
60
02
4a
01
24
c0
6a
02
69
fc
38
1a
00
ee
6a
00
69
fe
00
ee
4a
02
17
9e
48
2e
17
9a
00
ee
6a
01
00
ee
6a
00
69
fe
00
ee
4a
02
00
ee
60
04
49
fe
60
02
89
00
48
2e
69
00
49
04
6a
00
00
ee
60
00
4c
00
60
20
8c
00
67
04
00
ee
60
40
4c
40
60
60
8c
00
46
00
00
ee
67
fc
00
ee
60
01
f0
75
60
02
24
c0
24
c6
60
04
24
c0
24
c6
60
08
24
c0
60
1e
24
c6
00
e0
00
fd
00
00
00
00
00
00
00
00
00
00
00
00
00
00
00
00
00
00
00
00
00
00
00
00
00
00
00
00
00
00
00
00
2a
04
26
04
22
04
1e
04
1a
04
16
08
2e
fe
16
08
1a
04
1e
04
22
04
26
04
2a
10
2a
fd
22
03
22
ff
22
08
26
10
2e
fe
26
04
2a
04
2a
ff
2a
06
2a
ff
2a
06
26
0a
26
06
2e
fe
26
04
22
04
1e
03
1e
fd
1a
04
16
08
1a
ff
32
fe
2a
06
2a
1c
26
04
26
fc
1e
04
2e
fe
1a
05
16
04
2e
fe
26
08
26
ff
26
ff
1a
04
16
08
16
fd
2e
0e
16
08
2e
fe
16
04
2e
fe
16
03
2e
fe
16
04
16
fd
2e
fe
26
08
2e
06
2a
04
26
04
22
04
1e
04
1a
04
16
04
32
ff
32
ff
32
ff
32
ff
2e
08
1e
04
22
04
26
04
2a
04
32
fe
2e
04
2e
fd
2a
04
16
03
2a
1c
26
04
26
fb
32
fe
2a
04
26
04
22
04
1e
04
1a
04
16
04
1a
ff
22
ff
2a
ff
26
04
1e
04
32
fe
16
03
32
fe
1e
03
32
fe
16
03
16
fd
32
fe
1e
03
32
fe
16
03
2e
ff
2e
ff
2e
ff
2e
08
2a
04
16
06
2e
04
2a
04
26
04
22
04
1e
04
1a
04
16
08
16
fa
2e
04
2e
fd
22
03
1e
04
2e
02
26
02
16
03
1a
02
26
05
26
ff
2e
06
1a
03
1e
03
22
06
26
04
26
fd
16
06
32
fe
32
ff
2e
06
1a
03
16
03
1e
02
22
02
26
06
1a
04
1e
06
1e
fd
32
fe
26
04
16
03
22
03
1a
05
1a
ff
16
03
16
fd
2e
06
1e
02
1a
02
16
04
32
fe
1e
04
1e
fd
2e
08
2e
ff
2a
06
16
04
1a
01
16
01
1a
01
16
01
1a
01
16
01
1a
01
16
01
1a
01
16
01
1a
01
16
01
1a
01
16
01
1a
01
16
01
1a
01
16
01
1a
01
16
01
1a
01
16
01
1a
01
16
04
1a
04
1a
fd
16
04
32
fe
32
ff
2e
05
2a
02
26
03
22
02
1e
03
1a
02
16
03
1a
02
1e
ff
2e
06
22
02
16
08
16
fd
2e
06
16
03
2e
06
16
03
2e
06
16
03
2e
06
16
03
16
ff
16
02
2e
06
16
03
1e
fe
1a
05
1e
04
22
03
26
02
2a
01
2e
05
2e
ff
2a
04
2e
04
2e
ff
22
04
2e
05
2a
ff
2e
06
2e
ff
2e
05
2e
ff
2e
05
2e
ff
2a
04
32
fe
2e
03
2e
fd
2e
ff
1a
04
1e
fe
1a
04
2e
22
2e
f9
00
00
fe
00
00
00
00
00
00
00
68
27
20
64
1d
40
60
15
60
5c
0f
80
58
11
a0
54
0f
c0
50
15
e0
4c
1d
40
48
27
20
48
27
00
48
27
20
4c
1d
40
50
15
e0
54
0f
c0
58
11
a0
5c
0f
80
60
15
60
64
1d
40
68
27
20
68
27
00
00
0a
08
06
04
08
02
0a
08
00
06
08
0a
00
02
08
04
02
0a
08
00
11
00
0a
78
0e
dd
db
bf
ff
ff
ee
7a
e0
a5
50
a5
50
00
00
00
00
00
00
00
00
00
00
00
00
00
00
00
11
00
0a
78
0e
dd
db
bf
ff
ff
ee
39
f0
52
a8
52
a8
00
00
00
00
00
00
00
00
00
00
00
00
00
00
88
00
50
00
70
1e
db
bb
ff
fd
77
ff
07
5e
0a
a5
0a
a5
00
00
00
00
00
00
00
00
00
00
00
00
00
00
88
00
50
00
70
1e
db
bb
ff
fd
77
ff
0f
9c
15
4a
15
4a
00
00
00
00
00
00
00
00
00
00
00
00
00
00
f0
00
f0
50
e0
b0
e0
b0
f0
20
80
f0
f0
90
90
f0
00
80
00
c0
00
e0
00
f0
ff
f8
ff
fc
ff
fe
ff
ff
ff
fe
ff
fc
ff
f8
00
f0
00
e0
00
c0
00
80
00
00
f0
80
b0
a0
b0
a0
80
80
f0
00
10
a0
30
a0
00
00
f0
00
20
a0
a0
a0
00
00
f0
10
d0
b0
b0
d0
10
10
20
30
70
f0
00
00
00
00
00
00
00
00
00
1f
00
21
00
31
00
c1
03
2d
7c
8d
82
01
ff
ff
7f
ff
00
00
00
00
00
00
19
c0
26
20
40
10
80
08
81
08
40
88
20
44
20
42
40
42
80
82
80
02
40
0c
20
70
10
80
0f
00
00
00
00
00
01
e0
02
10
1c
10
20
08
40
08
83
88
84
44
88
02
40
02
40
02
80
02
80
04
43
08
24
90
18
60
00
00
00
f0
01
08
0e
04
30
02
40
01
41
01
42
02
42
04
22
04
11
02
10
81
10
01
08
02
04
64
03
98
06
18
09
24
10
c2
20
01
40
01
40
02
40
02
40
11
22
21
11
c1
10
02
10
04
08
38
08
40
07
80
00
00
01
f0
02
08
02
88
76
08
f2
08
59
f0
54
40
53
c0
70
60
00
50
00
48
00
a4
01
20
0a
10
04
08
00
10
00
00
00
00
03
e0
04
10
05
10
0c
10
04
10
3b
e0
78
80
2f
c0
28
a0
28
90
3b
90
02
80
02
e0
06
20
01
f0
02
08
02
88
76
08
f2
08
59
f2
54
44
53
f8
70
40
00
40
00
40
00
a0
01
10
0a
08
04
04
00
08
04
00
0a
00
11
20
20
a0
49
20
22
40
15
80
19
80
42
40
fc
20
50
1f
a8
11
14
10
08
10
00
30
00
00
00
00
04
00
02
02
79
05
85
08
85
10
87
e0
a5
10
85
08
79
04
12
02
04
04
1f
80
18
80
1f
80
08
00
10
00
20
20
10
50
08
80
05
00
02
00
02
00
02
0e
1f
ca
22
2a
4f
9a
10
4f
10
6e
11
40
10
40
0f
80
00
10
01
f8
01
18
01
f8
20
20
40
48
20
9e
10
a1
08
a5
07
e1
08
a1
10
a1
a0
9e
40
40
00
20
00
00
14
00
0e
20
14
50
2d
88
55
24
24
82
02
44
01
a8
01
90
02
40
84
38
f8
00
08
00
08
00
08
00
18
00
0f
80
10
40
11
40
10
6e
10
4f
0f
9a
02
2a
07
ca
0a
0e
12
00
12
00
05
00
08
80
10
50
20
20
10
00
0f
80
10
40
11
40
10
6e
10
4f
0f
9a
02
2a
07
ca
06
0e
06
00
03
00
02
00
02
00
06
00
0a
00
07
00
01
f0
02
08
02
88
76
08
f2
08
59
f0
54
40
53
e0
70
50
00
48
00
48
00
a0
01
10
0a
08
04
04
00
08
01
f0
02
08
02
88
76
08
f2
08
59
f0
54
40
53
e0
70
60
00
60
00
c0
00
40
00
40
00
60
00
50
00
e0
3c
00
6b
00
d5
40
aa
a8
d5
55
aa
a8
d5
40
6b
00
3c
00
00
00
00
00
00
00
00
00
00
00
00
00
00
00
00
00
07
c0
18
30
20
08
40
04
4c
64
9e
f2
96
b2
8c
62
80
02
80
02
43
84
44
44
20
08
18
30
07
c0
00
00
07
c0
18
30
20
08
40
c4
41
e4
81
a2
8c
c2
9e
02
9a
1a
8c
22
40
44
40
84
20
88
18
30
07
c0
00
00
07
c0
18
30
20
08
46
04
4f
04
8d
12
86
22
80
22
86
22
8f
12
4d
04
46
04
20
08
18
30
07
c0
00
00
07
c0
18
30
20
88
40
84
4c
44
9a
22
9e
1a
8c
02
81
82
83
42
43
c4
41
84
20
08
18
30
07
c0
00
00
07
c0
18
30
20
08
44
44
43
84
80
02
80
02
8c
62
9a
d2
9e
f2
4c
64
40
04
20
08
18
30
07
c0
00
00
07
c0
18
30
22
08
42
04
44
64
88
b2
b0
f2
80
62
83
02
85
82
47
84
43
04
20
08
18
30
07
c0
00
00
07
c0
18
30
20
08
40
c4
41
64
91
e2
88
c2
88
02
88
c2
91
62
41
e4
40
c4
20
08
18
30
07
c0
00
00
07
c0
18
30
20
08
43
04
47
84
85
82
83
02
80
62
b0
f2
88
b2
44
64
42
04
22
08
18
30
07
c0
