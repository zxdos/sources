-- ZPU
--
-- Copyright 2004-2008 oharboe - �yvind Harboe - oyvind.harboe@zylin.com
-- Modified by Alastair M. Robinson for the ZPUFlex project.
--
-- The FreeBSD license
-- 
-- Redistribution and use in source and binary forms, with or without
-- modification, are permitted provided that the following conditions
-- are met:
-- 
-- 1. Redistributions of source code must retain the above copyright
--    notice, this list of conditions and the following disclaimer.
-- 2. Redistributions in binary form must reproduce the above
--    copyright notice, this list of conditions and the following
--    disclaimer in the documentation and/or other materials
--    provided with the distribution.
-- 
-- THIS SOFTWARE IS PROVIDED BY THE ZPU PROJECT ``AS IS'' AND ANY
-- EXPRESS OR IMPLIED WARRANTIES, INCLUDING, BUT NOT LIMITED TO,
-- THE IMPLIED WARRANTIES OF MERCHANTABILITY AND FITNESS FOR A
-- PARTICULAR PURPOSE ARE DISCLAIMED. IN NO EVENT SHALL THE
-- ZPU PROJECT OR CONTRIBUTORS BE LIABLE FOR ANY DIRECT,
-- INDIRECT, INCIDENTAL, SPECIAL, EXEMPLARY, OR CONSEQUENTIAL DAMAGES
-- (INCLUDING, BUT NOT LIMITED TO, PROCUREMENT OF SUBSTITUTE GOODS
-- OR SERVICES; LOSS OF USE, DATA, OR PROFITS; OR BUSINESS INTERRUPTION)
-- HOWEVER CAUSED AND ON ANY THEORY OF LIABILITY, WHETHER IN CONTRACT,
-- STRICT LIABILITY, OR TORT (INCLUDING NEGLIGENCE OR OTHERWISE)
-- ARISING IN ANY WAY OUT OF THE USE OF THIS SOFTWARE, EVEN IF
-- ADVISED OF THE POSSIBILITY OF SUCH DAMAGE.
-- 
-- The views and conclusions contained in the software and documentation
-- are those of the authors and should not be interpreted as representing
-- official policies, either expressed or implied, of the ZPU Project.

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;


library work;
use work.zpupkg.all;

entity CtrlROM_ROM is
generic
	(
		maxAddrBitBRAM : integer := maxAddrBitBRAMLimit -- Specify your actual ROM size to save LEs and unnecessary block RAM usage.
	);
port (
	clk : in std_logic;
	areset : in std_logic := '0';
	from_zpu : in ZPU_ToROM;
	to_zpu : out ZPU_FromROM
);
end CtrlROM_ROM;

architecture arch of CtrlROM_ROM is

type ram_type is array(natural range 0 to ((2**(maxAddrBitBRAM+1))/4)-1) of std_logic_vector(wordSize-1 downto 0);

shared variable ram : ram_type :=
(
     0 => x"0b0b0b0b",
     1 => x"8c0b0b0b",
     2 => x"0b81e004",
     3 => x"0b0b0b0b",
     4 => x"8c04ff0d",
     5 => x"80040400",
     6 => x"00000016",
     7 => x"00000000",
     8 => x"0b0b80c8",
     9 => x"d4080b0b",
    10 => x"80c8d808",
    11 => x"0b0b80c8",
    12 => x"dc080b0b",
    13 => x"0b0b9808",
    14 => x"2d0b0b80",
    15 => x"c8dc0c0b",
    16 => x"0b80c8d8",
    17 => x"0c0b0b80",
    18 => x"c8d40c04",
    19 => x"00000000",
    20 => x"00000000",
    21 => x"00000000",
    22 => x"00000000",
    23 => x"00000000",
    24 => x"71fd0608",
    25 => x"72830609",
    26 => x"81058205",
    27 => x"832b2a83",
    28 => x"ffff0652",
    29 => x"0471fc06",
    30 => x"08728306",
    31 => x"09810583",
    32 => x"05101010",
    33 => x"2a81ff06",
    34 => x"520471fd",
    35 => x"060883ff",
    36 => x"ff738306",
    37 => x"09810582",
    38 => x"05832b2b",
    39 => x"09067383",
    40 => x"ffff0673",
    41 => x"83060981",
    42 => x"05820583",
    43 => x"2b0b2b07",
    44 => x"72fc060c",
    45 => x"51510471",
    46 => x"fc06080b",
    47 => x"0b0bbaa8",
    48 => x"73830610",
    49 => x"10050806",
    50 => x"7381ff06",
    51 => x"73830609",
    52 => x"81058305",
    53 => x"1010102b",
    54 => x"0772fc06",
    55 => x"0c515104",
    56 => x"80c8d470",
    57 => x"80d69c27",
    58 => x"8b388071",
    59 => x"70840553",
    60 => x"0c81e304",
    61 => x"8c5189f5",
    62 => x"0402fc05",
    63 => x"0df88051",
    64 => x"8f0b80c8",
    65 => x"e40c9f0b",
    66 => x"80c8e80c",
    67 => x"a0717081",
    68 => x"05533480",
    69 => x"c8e808ff",
    70 => x"0580c8e8",
    71 => x"0c80c8e8",
    72 => x"088025e8",
    73 => x"3880c8e4",
    74 => x"08ff0580",
    75 => x"c8e40c80",
    76 => x"c8e40880",
    77 => x"25d03880",
    78 => x"0b80c8e8",
    79 => x"0c800b80",
    80 => x"c8e40c02",
    81 => x"84050d04",
    82 => x"02f0050d",
    83 => x"f88053f8",
    84 => x"a05483bf",
    85 => x"52737081",
    86 => x"05553351",
    87 => x"70737081",
    88 => x"055534ff",
    89 => x"12527180",
    90 => x"25eb38fb",
    91 => x"c0539f52",
    92 => x"a0737081",
    93 => x"055534ff",
    94 => x"12527180",
    95 => x"25f23802",
    96 => x"90050d04",
    97 => x"02f4050d",
    98 => x"74538e0b",
    99 => x"80c8e408",
   100 => x"25913882",
   101 => x"c82d80c8",
   102 => x"e408ff05",
   103 => x"80c8e40c",
   104 => x"838a0480",
   105 => x"c8e40880",
   106 => x"c8e80853",
   107 => x"51728a2e",
   108 => x"098106be",
   109 => x"38715171",
   110 => x"9f24a438",
   111 => x"80c8e408",
   112 => x"a02911f8",
   113 => x"80115151",
   114 => x"a0713480",
   115 => x"c8e80881",
   116 => x"0580c8e8",
   117 => x"0c80c8e8",
   118 => x"08519f71",
   119 => x"25de3880",
   120 => x"0b80c8e8",
   121 => x"0c80c8e4",
   122 => x"08810580",
   123 => x"c8e40c84",
   124 => x"880470a0",
   125 => x"2912f880",
   126 => x"11515172",
   127 => x"713480c8",
   128 => x"e8088105",
   129 => x"80c8e80c",
   130 => x"80c8e808",
   131 => x"a02e0981",
   132 => x"06913880",
   133 => x"0b80c8e8",
   134 => x"0c80c8e4",
   135 => x"08810580",
   136 => x"c8e40c02",
   137 => x"8c050d04",
   138 => x"02e8050d",
   139 => x"77795656",
   140 => x"880bfc16",
   141 => x"77712c8f",
   142 => x"06545254",
   143 => x"80537272",
   144 => x"25953871",
   145 => x"53fbe014",
   146 => x"51877134",
   147 => x"8114ff14",
   148 => x"545472f1",
   149 => x"387153f9",
   150 => x"1576712c",
   151 => x"87065351",
   152 => x"71802e8b",
   153 => x"38fbe014",
   154 => x"51717134",
   155 => x"81145472",
   156 => x"8e249538",
   157 => x"8f733153",
   158 => x"fbe01451",
   159 => x"a0713481",
   160 => x"14ff1454",
   161 => x"5472f138",
   162 => x"0298050d",
   163 => x"0402ec05",
   164 => x"0d800b80",
   165 => x"c8ec0cf6",
   166 => x"8c08f690",
   167 => x"0871882c",
   168 => x"555381ff",
   169 => x"06547274",
   170 => x"25893873",
   171 => x"53820b80",
   172 => x"c8ec0c71",
   173 => x"882c7281",
   174 => x"ff065355",
   175 => x"7472258d",
   176 => x"387180c8",
   177 => x"ec088407",
   178 => x"80c8ec0c",
   179 => x"5572842b",
   180 => x"75832b56",
   181 => x"5386a073",
   182 => x"258f3883",
   183 => x"0b0b0b80",
   184 => x"c18c0c80",
   185 => x"e35485f4",
   186 => x"04810b0b",
   187 => x"0b80c18c",
   188 => x"0c828554",
   189 => x"810b0b0b",
   190 => x"80c18c08",
   191 => x"2bff05f6",
   192 => x"880cfc08",
   193 => x"ff941670",
   194 => x"9f2a1170",
   195 => x"812c80c8",
   196 => x"ec085255",
   197 => x"51515176",
   198 => x"802e8538",
   199 => x"70810751",
   200 => x"70f6940c",
   201 => x"73098105",
   202 => x"f6800c71",
   203 => x"098105f6",
   204 => x"840c0294",
   205 => x"050d0402",
   206 => x"f4050d74",
   207 => x"53727081",
   208 => x"055480f5",
   209 => x"2d527180",
   210 => x"2e893871",
   211 => x"5183842d",
   212 => x"86bd0481",
   213 => x"0b80c8d4",
   214 => x"0c028c05",
   215 => x"0d0402fc",
   216 => x"050d8180",
   217 => x"8051c011",
   218 => x"5170fb38",
   219 => x"0284050d",
   220 => x"0402fc05",
   221 => x"0dec5183",
   222 => x"710c86de",
   223 => x"2d82710c",
   224 => x"0284050d",
   225 => x"0402fc05",
   226 => x"0d84bf51",
   227 => x"86de2dff",
   228 => x"11517080",
   229 => x"25f63802",
   230 => x"84050d04",
   231 => x"0402fc05",
   232 => x"0d8fe32d",
   233 => x"80c8d408",
   234 => x"80c6900c",
   235 => x"80c4f851",
   236 => x"92982d02",
   237 => x"84050d04",
   238 => x"02fc050d",
   239 => x"8fe32d80",
   240 => x"c8d40880",
   241 => x"c4e80c80",
   242 => x"c3d05192",
   243 => x"982d0284",
   244 => x"050d0402",
   245 => x"dc050d7a",
   246 => x"54805984",
   247 => x"0bec0c80",
   248 => x"c8fc0882",
   249 => x"80078280",
   250 => x"327080c8",
   251 => x"fc0cfc0c",
   252 => x"86de2d73",
   253 => x"5280c8f0",
   254 => x"51b18d2d",
   255 => x"80c8d408",
   256 => x"792e81ac",
   257 => x"3880c8f4",
   258 => x"08557485",
   259 => x"2e098106",
   260 => x"a5387351",
   261 => x"86b72d87",
   262 => x"852d8785",
   263 => x"2d87852d",
   264 => x"87852d87",
   265 => x"852d8785",
   266 => x"2d80cc88",
   267 => x"08519298",
   268 => x"2d815389",
   269 => x"eb0474f8",
   270 => x"0ca50bec",
   271 => x"0c87852d",
   272 => x"840bec0c",
   273 => x"78ff1655",
   274 => x"5873802e",
   275 => x"8b388118",
   276 => x"74812a55",
   277 => x"5888c904",
   278 => x"f7185881",
   279 => x"59807525",
   280 => x"80ce3877",
   281 => x"52735184",
   282 => x"a82d80cc",
   283 => x"d45280c8",
   284 => x"f051b3da",
   285 => x"2d80c8d4",
   286 => x"08802e9b",
   287 => x"3880ccd4",
   288 => x"5783fc56",
   289 => x"76708405",
   290 => x"5808e80c",
   291 => x"fc165675",
   292 => x"8025f138",
   293 => x"899f0480",
   294 => x"c8d40859",
   295 => x"84805580",
   296 => x"c8f051b3",
   297 => x"aa2dfc80",
   298 => x"15811555",
   299 => x"5588dd04",
   300 => x"800b80c1",
   301 => x"900c80c8",
   302 => x"fc088280",
   303 => x"07828032",
   304 => x"7080c8fc",
   305 => x"0cfc0c78",
   306 => x"802e9738",
   307 => x"80cc8808",
   308 => x"5192982d",
   309 => x"810bec0c",
   310 => x"87852d82",
   311 => x"0bec0c89",
   312 => x"e90480c3",
   313 => x"ac519298",
   314 => x"2d785372",
   315 => x"80c8d40c",
   316 => x"02a4050d",
   317 => x"0402f405",
   318 => x"0d840b80",
   319 => x"c8fc0c80",
   320 => x"5186f12d",
   321 => x"840bec0c",
   322 => x"8fb32d8b",
   323 => x"de2d81f9",
   324 => x"2d83528f",
   325 => x"962d8151",
   326 => x"858d2dff",
   327 => x"12527180",
   328 => x"25f13884",
   329 => x"0bec0cbf",
   330 => x"c05186b7",
   331 => x"2da7c52d",
   332 => x"80c8d408",
   333 => x"802e818f",
   334 => x"38810bec",
   335 => x"0c840bec",
   336 => x"0c87d351",
   337 => x"baa22d80",
   338 => x"c8fc0870",
   339 => x"822c80c6",
   340 => x"e80cfc0c",
   341 => x"80ccb408",
   342 => x"882a7081",
   343 => x"06515271",
   344 => x"802e8c38",
   345 => x"80c2c00b",
   346 => x"80cc880c",
   347 => x"8af70480",
   348 => x"c1940b80",
   349 => x"cc880c80",
   350 => x"cc880851",
   351 => x"92982d84",
   352 => x"0b80ccc8",
   353 => x"0c8fec2d",
   354 => x"8bea2d92",
   355 => x"ab2d80cc",
   356 => x"8808ac11",
   357 => x"80f52d70",
   358 => x"80c8fc0c",
   359 => x"80c6e808",
   360 => x"81065254",
   361 => x"5271802e",
   362 => x"88387284",
   363 => x"0780c8fc",
   364 => x"0c80c8fc",
   365 => x"08fc0c86",
   366 => x"5280c8d4",
   367 => x"08833884",
   368 => x"5271ec0c",
   369 => x"8b880480",
   370 => x"0b80c8d4",
   371 => x"0c028c05",
   372 => x"0d047198",
   373 => x"0c04ffb0",
   374 => x"0880c8d4",
   375 => x"0c04810b",
   376 => x"ffb00c04",
   377 => x"800bffb0",
   378 => x"0c0402f4",
   379 => x"050d8cf8",
   380 => x"0480c8d4",
   381 => x"0881f02e",
   382 => x"0981068a",
   383 => x"38810b80",
   384 => x"c6e00c8c",
   385 => x"f80480c8",
   386 => x"d40881e0",
   387 => x"2e098106",
   388 => x"8a38810b",
   389 => x"80c6e40c",
   390 => x"8cf80480",
   391 => x"c8d40852",
   392 => x"80c6e408",
   393 => x"802e8938",
   394 => x"80c8d408",
   395 => x"81800552",
   396 => x"71842c72",
   397 => x"8f065353",
   398 => x"80c6e008",
   399 => x"802e9a38",
   400 => x"72842980",
   401 => x"c6a00572",
   402 => x"1381712b",
   403 => x"70097308",
   404 => x"06730c51",
   405 => x"53538cec",
   406 => x"04728429",
   407 => x"80c6a005",
   408 => x"72138371",
   409 => x"2b720807",
   410 => x"720c5353",
   411 => x"800b80c6",
   412 => x"e40c800b",
   413 => x"80c6e00c",
   414 => x"80cc8c51",
   415 => x"8dff2d80",
   416 => x"c8d408ff",
   417 => x"24feea38",
   418 => x"800b80c8",
   419 => x"d40c028c",
   420 => x"050d0402",
   421 => x"f8050d80",
   422 => x"c6a0528f",
   423 => x"51807270",
   424 => x"8405540c",
   425 => x"ff115170",
   426 => x"8025f238",
   427 => x"0288050d",
   428 => x"0402f005",
   429 => x"0d75518b",
   430 => x"e42d7082",
   431 => x"2cfc0680",
   432 => x"c6a01172",
   433 => x"109e0671",
   434 => x"0870722a",
   435 => x"70830682",
   436 => x"742b7009",
   437 => x"7406760c",
   438 => x"54515657",
   439 => x"5351538b",
   440 => x"de2d7180",
   441 => x"c8d40c02",
   442 => x"90050d04",
   443 => x"02fc050d",
   444 => x"72518071",
   445 => x"0c800b84",
   446 => x"120c0284",
   447 => x"050d0402",
   448 => x"f0050d75",
   449 => x"70088412",
   450 => x"08535353",
   451 => x"ff547171",
   452 => x"2ea8388b",
   453 => x"e42d8413",
   454 => x"08708429",
   455 => x"14881170",
   456 => x"087081ff",
   457 => x"06841808",
   458 => x"81118706",
   459 => x"841a0c53",
   460 => x"51555151",
   461 => x"518bde2d",
   462 => x"71547380",
   463 => x"c8d40c02",
   464 => x"90050d04",
   465 => x"02f4050d",
   466 => x"8be42de0",
   467 => x"08708b2a",
   468 => x"70810651",
   469 => x"52537080",
   470 => x"2ea13880",
   471 => x"cc8c0870",
   472 => x"842980cc",
   473 => x"94057481",
   474 => x"ff06710c",
   475 => x"515180cc",
   476 => x"8c088111",
   477 => x"870680cc",
   478 => x"8c0c5172",
   479 => x"8c2c83ff",
   480 => x"0680ccb4",
   481 => x"0c800b80",
   482 => x"ccb80c8b",
   483 => x"d62d8bde",
   484 => x"2d028c05",
   485 => x"0d0402fc",
   486 => x"050d8be4",
   487 => x"2d810b80",
   488 => x"ccb80c8b",
   489 => x"de2d80cc",
   490 => x"b8085170",
   491 => x"f9380284",
   492 => x"050d0402",
   493 => x"fc050d80",
   494 => x"cc8c518d",
   495 => x"ec2d8d93",
   496 => x"2d8ec451",
   497 => x"8bd22d02",
   498 => x"84050d04",
   499 => x"02fc050d",
   500 => x"8fcf5186",
   501 => x"de2dff11",
   502 => x"51708025",
   503 => x"f6380284",
   504 => x"050d0480",
   505 => x"ccc00880",
   506 => x"c8d40c04",
   507 => x"02fc050d",
   508 => x"810b80c7",
   509 => x"940c8151",
   510 => x"858d2d02",
   511 => x"84050d04",
   512 => x"02fc050d",
   513 => x"908a048b",
   514 => x"ea2d80f6",
   515 => x"518db12d",
   516 => x"80c8d408",
   517 => x"f23880da",
   518 => x"518db12d",
   519 => x"80c8d408",
   520 => x"e63880c7",
   521 => x"9008518d",
   522 => x"b12d80c8",
   523 => x"d408d838",
   524 => x"80c8d408",
   525 => x"80c7940c",
   526 => x"80c8d408",
   527 => x"51858d2d",
   528 => x"0284050d",
   529 => x"0402ec05",
   530 => x"0d765480",
   531 => x"52870b88",
   532 => x"1580f52d",
   533 => x"56537472",
   534 => x"248338a0",
   535 => x"53725183",
   536 => x"842d8112",
   537 => x"8b1580f5",
   538 => x"2d545272",
   539 => x"7225de38",
   540 => x"0294050d",
   541 => x"0402f005",
   542 => x"0d80ccc0",
   543 => x"085481f9",
   544 => x"2d800b80",
   545 => x"ccc40c73",
   546 => x"08802e81",
   547 => x"8638820b",
   548 => x"80c8e80c",
   549 => x"80ccc408",
   550 => x"8f0680c8",
   551 => x"e40c7308",
   552 => x"5271832e",
   553 => x"96387183",
   554 => x"26893871",
   555 => x"812eaf38",
   556 => x"91fc0471",
   557 => x"852e9f38",
   558 => x"91fc0488",
   559 => x"1480f52d",
   560 => x"841508bf",
   561 => x"d8535452",
   562 => x"86b72d71",
   563 => x"84291370",
   564 => x"08525292",
   565 => x"80047351",
   566 => x"90c52d91",
   567 => x"fc0480c6",
   568 => x"e8088815",
   569 => x"082c7081",
   570 => x"06515271",
   571 => x"802e8738",
   572 => x"bfdc5191",
   573 => x"f904bfe0",
   574 => x"5186b72d",
   575 => x"84140851",
   576 => x"86b72d80",
   577 => x"ccc40881",
   578 => x"0580ccc4",
   579 => x"0c8c1454",
   580 => x"91870402",
   581 => x"90050d04",
   582 => x"7180ccc0",
   583 => x"0c90f52d",
   584 => x"80ccc408",
   585 => x"ff0580cc",
   586 => x"c80c0402",
   587 => x"e8050d80",
   588 => x"ccc00880",
   589 => x"cccc0857",
   590 => x"5580f651",
   591 => x"8db12d80",
   592 => x"c8d40881",
   593 => x"2a708106",
   594 => x"51527180",
   595 => x"2ea23892",
   596 => x"d5048bea",
   597 => x"2d80f651",
   598 => x"8db12d80",
   599 => x"c8d408f2",
   600 => x"3880c794",
   601 => x"08813270",
   602 => x"80c7940c",
   603 => x"51858d2d",
   604 => x"800b80cc",
   605 => x"bc0c8651",
   606 => x"8db12d80",
   607 => x"c8d40881",
   608 => x"2a708106",
   609 => x"51527180",
   610 => x"2e8b3880",
   611 => x"c8fc0890",
   612 => x"3280c8fc",
   613 => x"0c8c518d",
   614 => x"b12d80c8",
   615 => x"d408812a",
   616 => x"70810651",
   617 => x"5271802e",
   618 => x"80d13880",
   619 => x"c6ec0880",
   620 => x"c7800880",
   621 => x"c6ec0c80",
   622 => x"c7800c80",
   623 => x"c6f00880",
   624 => x"c7840880",
   625 => x"c6f00c80",
   626 => x"c7840c80",
   627 => x"c6f40880",
   628 => x"c7880880",
   629 => x"c6f40c80",
   630 => x"c7880c80",
   631 => x"c6f80880",
   632 => x"c78c0880",
   633 => x"c6f80c80",
   634 => x"c78c0c80",
   635 => x"c6fc0880",
   636 => x"c7900880",
   637 => x"c6fc0c80",
   638 => x"c7900c80",
   639 => x"ccb408a0",
   640 => x"06528072",
   641 => x"2596388f",
   642 => x"cc2d8bea",
   643 => x"2d80c794",
   644 => x"08813270",
   645 => x"80c7940c",
   646 => x"51858d2d",
   647 => x"80c79408",
   648 => x"82ef3880",
   649 => x"c7800851",
   650 => x"8db12d80",
   651 => x"c8d40880",
   652 => x"2e8b3880",
   653 => x"ccbc0881",
   654 => x"0780ccbc",
   655 => x"0c80c784",
   656 => x"08518db1",
   657 => x"2d80c8d4",
   658 => x"08802e8b",
   659 => x"3880ccbc",
   660 => x"08820780",
   661 => x"ccbc0c80",
   662 => x"c7880851",
   663 => x"8db12d80",
   664 => x"c8d40880",
   665 => x"2e8b3880",
   666 => x"ccbc0884",
   667 => x"0780ccbc",
   668 => x"0c80c78c",
   669 => x"08518db1",
   670 => x"2d80c8d4",
   671 => x"08802e8b",
   672 => x"3880ccbc",
   673 => x"08880780",
   674 => x"ccbc0c80",
   675 => x"c7900851",
   676 => x"8db12d80",
   677 => x"c8d40880",
   678 => x"2e8b3880",
   679 => x"ccbc0890",
   680 => x"0780ccbc",
   681 => x"0c80c6ec",
   682 => x"08518db1",
   683 => x"2d80c8d4",
   684 => x"08802e8c",
   685 => x"3880ccbc",
   686 => x"08828007",
   687 => x"80ccbc0c",
   688 => x"80c6f008",
   689 => x"518db12d",
   690 => x"80c8d408",
   691 => x"802e8c38",
   692 => x"80ccbc08",
   693 => x"84800780",
   694 => x"ccbc0c80",
   695 => x"c6f40851",
   696 => x"8db12d80",
   697 => x"c8d40880",
   698 => x"2e8c3880",
   699 => x"ccbc0888",
   700 => x"800780cc",
   701 => x"bc0c80c6",
   702 => x"f808518d",
   703 => x"b12d80c8",
   704 => x"d408802e",
   705 => x"8c3880cc",
   706 => x"bc089080",
   707 => x"0780ccbc",
   708 => x"0c80c6fc",
   709 => x"08518db1",
   710 => x"2d80c8d4",
   711 => x"08802e8c",
   712 => x"3880ccbc",
   713 => x"08a08007",
   714 => x"80ccbc0c",
   715 => x"94518db1",
   716 => x"2d80c8d4",
   717 => x"08529151",
   718 => x"8db12d71",
   719 => x"80c8d408",
   720 => x"065280e6",
   721 => x"518db12d",
   722 => x"7180c8d4",
   723 => x"08065271",
   724 => x"802e8d38",
   725 => x"80ccbc08",
   726 => x"84808007",
   727 => x"80ccbc0c",
   728 => x"80fe518d",
   729 => x"b12d80c8",
   730 => x"d4085287",
   731 => x"518db12d",
   732 => x"7180c8d4",
   733 => x"08075271",
   734 => x"802e8d38",
   735 => x"80ccbc08",
   736 => x"88808007",
   737 => x"80ccbc0c",
   738 => x"80ccbc08",
   739 => x"ed0c9f9c",
   740 => x"0494518d",
   741 => x"b12d80c8",
   742 => x"d4085291",
   743 => x"518db12d",
   744 => x"7180c8d4",
   745 => x"08065280",
   746 => x"e6518db1",
   747 => x"2d7180c8",
   748 => x"d4080652",
   749 => x"71802e8d",
   750 => x"3880ccbc",
   751 => x"08848080",
   752 => x"0780ccbc",
   753 => x"0c80fe51",
   754 => x"8db12d80",
   755 => x"c8d40852",
   756 => x"87518db1",
   757 => x"2d7180c8",
   758 => x"d4080752",
   759 => x"71802e8d",
   760 => x"3880ccbc",
   761 => x"08888080",
   762 => x"0780ccbc",
   763 => x"0c80ccbc",
   764 => x"08ed0c81",
   765 => x"f5518db1",
   766 => x"2d80c8d4",
   767 => x"08812a70",
   768 => x"81065152",
   769 => x"71a43880",
   770 => x"c7800851",
   771 => x"8db12d80",
   772 => x"c8d40881",
   773 => x"2a708106",
   774 => x"5152718e",
   775 => x"3880ccb4",
   776 => x"08810652",
   777 => x"80722580",
   778 => x"c23880cc",
   779 => x"b4088106",
   780 => x"52807225",
   781 => x"84388fcc",
   782 => x"2d80ccc8",
   783 => x"08527180",
   784 => x"2e8a38ff",
   785 => x"1280ccc8",
   786 => x"0c98eb04",
   787 => x"80ccc408",
   788 => x"1080ccc4",
   789 => x"08057084",
   790 => x"29165152",
   791 => x"88120880",
   792 => x"2e8938ff",
   793 => x"51881208",
   794 => x"52712d81",
   795 => x"f2518db1",
   796 => x"2d80c8d4",
   797 => x"08812a70",
   798 => x"81065152",
   799 => x"71a43880",
   800 => x"c7840851",
   801 => x"8db12d80",
   802 => x"c8d40881",
   803 => x"2a708106",
   804 => x"5152718e",
   805 => x"3880ccb4",
   806 => x"08820652",
   807 => x"80722580",
   808 => x"c33880cc",
   809 => x"b4088206",
   810 => x"52807225",
   811 => x"84388fcc",
   812 => x"2d80ccc4",
   813 => x"08ff1180",
   814 => x"ccc80856",
   815 => x"53537372",
   816 => x"258a3881",
   817 => x"1480ccc8",
   818 => x"0c99e404",
   819 => x"72101370",
   820 => x"84291651",
   821 => x"52881208",
   822 => x"802e8938",
   823 => x"fe518812",
   824 => x"0852712d",
   825 => x"81fd518d",
   826 => x"b12d80c8",
   827 => x"d408812a",
   828 => x"70810651",
   829 => x"5271a438",
   830 => x"80c78808",
   831 => x"518db12d",
   832 => x"80c8d408",
   833 => x"812a7081",
   834 => x"06515271",
   835 => x"8e3880cc",
   836 => x"b4088406",
   837 => x"52807225",
   838 => x"80c03880",
   839 => x"ccb40884",
   840 => x"06528072",
   841 => x"2584388f",
   842 => x"cc2d80cc",
   843 => x"c808802e",
   844 => x"8a38800b",
   845 => x"80ccc80c",
   846 => x"9ada0480",
   847 => x"ccc40810",
   848 => x"80ccc408",
   849 => x"05708429",
   850 => x"16515288",
   851 => x"1208802e",
   852 => x"8938fd51",
   853 => x"88120852",
   854 => x"712d81fa",
   855 => x"518db12d",
   856 => x"80c8d408",
   857 => x"812a7081",
   858 => x"06515271",
   859 => x"a43880c7",
   860 => x"8c08518d",
   861 => x"b12d80c8",
   862 => x"d408812a",
   863 => x"70810651",
   864 => x"52718e38",
   865 => x"80ccb408",
   866 => x"88065280",
   867 => x"722580c0",
   868 => x"3880ccb4",
   869 => x"08880652",
   870 => x"80722584",
   871 => x"388fcc2d",
   872 => x"80ccc408",
   873 => x"ff115452",
   874 => x"80ccc808",
   875 => x"73258938",
   876 => x"7280ccc8",
   877 => x"0c9bd004",
   878 => x"71101270",
   879 => x"84291651",
   880 => x"52881208",
   881 => x"802e8938",
   882 => x"fc518812",
   883 => x"0852712d",
   884 => x"80ccc808",
   885 => x"70535473",
   886 => x"802e8a38",
   887 => x"8c15ff15",
   888 => x"55559bd7",
   889 => x"04820b80",
   890 => x"c8e80c71",
   891 => x"8f0680c8",
   892 => x"e40c81eb",
   893 => x"518db12d",
   894 => x"80c8d408",
   895 => x"812a7081",
   896 => x"06515271",
   897 => x"802ead38",
   898 => x"7408852e",
   899 => x"098106a4",
   900 => x"38881580",
   901 => x"f52dff05",
   902 => x"52718816",
   903 => x"81b72d71",
   904 => x"982b5271",
   905 => x"80258838",
   906 => x"800b8816",
   907 => x"81b72d74",
   908 => x"5190c52d",
   909 => x"81f4518d",
   910 => x"b12d80c8",
   911 => x"d408812a",
   912 => x"70810651",
   913 => x"5271802e",
   914 => x"b3387408",
   915 => x"852e0981",
   916 => x"06aa3888",
   917 => x"1580f52d",
   918 => x"81055271",
   919 => x"881681b7",
   920 => x"2d7181ff",
   921 => x"068b1680",
   922 => x"f52d5452",
   923 => x"72722787",
   924 => x"38728816",
   925 => x"81b72d74",
   926 => x"5190c52d",
   927 => x"80da518d",
   928 => x"b12d80c8",
   929 => x"d408812a",
   930 => x"70810651",
   931 => x"52718e38",
   932 => x"80ccb408",
   933 => x"90065280",
   934 => x"722581bc",
   935 => x"3880ccc0",
   936 => x"0880ccb4",
   937 => x"08900653",
   938 => x"53807225",
   939 => x"84388fcc",
   940 => x"2d80ccc8",
   941 => x"08547380",
   942 => x"2e8a388c",
   943 => x"13ff1555",
   944 => x"539db604",
   945 => x"72085271",
   946 => x"822ea638",
   947 => x"71822689",
   948 => x"3871812e",
   949 => x"aa389ed8",
   950 => x"0471832e",
   951 => x"b4387184",
   952 => x"2e098106",
   953 => x"80f23888",
   954 => x"13085192",
   955 => x"982d9ed8",
   956 => x"0480ccc8",
   957 => x"08518813",
   958 => x"0852712d",
   959 => x"9ed80481",
   960 => x"0b881408",
   961 => x"2b80c6e8",
   962 => x"083280c6",
   963 => x"e80c9eac",
   964 => x"04881380",
   965 => x"f52d8105",
   966 => x"8b1480f5",
   967 => x"2d535471",
   968 => x"74248338",
   969 => x"80547388",
   970 => x"1481b72d",
   971 => x"90f52d9e",
   972 => x"d8047508",
   973 => x"802ea438",
   974 => x"7508518d",
   975 => x"b12d80c8",
   976 => x"d4088106",
   977 => x"5271802e",
   978 => x"8c3880cc",
   979 => x"c8085184",
   980 => x"16085271",
   981 => x"2d881656",
   982 => x"75d83880",
   983 => x"54800b80",
   984 => x"c8e80c73",
   985 => x"8f0680c8",
   986 => x"e40ca052",
   987 => x"7380ccc8",
   988 => x"082e0981",
   989 => x"06993880",
   990 => x"ccc408ff",
   991 => x"05743270",
   992 => x"09810570",
   993 => x"72079f2a",
   994 => x"91713151",
   995 => x"51535371",
   996 => x"5183842d",
   997 => x"8114548e",
   998 => x"7425c238",
   999 => x"80c79408",
  1000 => x"80c8d40c",
  1001 => x"0298050d",
  1002 => x"0402f405",
  1003 => x"0dd45281",
  1004 => x"ff720c71",
  1005 => x"085381ff",
  1006 => x"720c7288",
  1007 => x"2b83fe80",
  1008 => x"06720870",
  1009 => x"81ff0651",
  1010 => x"525381ff",
  1011 => x"720c7271",
  1012 => x"07882b72",
  1013 => x"087081ff",
  1014 => x"06515253",
  1015 => x"81ff720c",
  1016 => x"72710788",
  1017 => x"2b720870",
  1018 => x"81ff0672",
  1019 => x"0780c8d4",
  1020 => x"0c525302",
  1021 => x"8c050d04",
  1022 => x"02f4050d",
  1023 => x"74767181",
  1024 => x"ff06d40c",
  1025 => x"535380cc",
  1026 => x"d0088538",
  1027 => x"71892b52",
  1028 => x"71982ad4",
  1029 => x"0c71902a",
  1030 => x"7081ff06",
  1031 => x"d40c5171",
  1032 => x"882a7081",
  1033 => x"ff06d40c",
  1034 => x"517181ff",
  1035 => x"06d40c72",
  1036 => x"902a7081",
  1037 => x"ff06d40c",
  1038 => x"51d40870",
  1039 => x"81ff0651",
  1040 => x"5182b8bf",
  1041 => x"527081ff",
  1042 => x"2e098106",
  1043 => x"943881ff",
  1044 => x"0bd40cd4",
  1045 => x"087081ff",
  1046 => x"06ff1454",
  1047 => x"515171e5",
  1048 => x"387080c8",
  1049 => x"d40c028c",
  1050 => x"050d0402",
  1051 => x"fc050d81",
  1052 => x"c75181ff",
  1053 => x"0bd40cff",
  1054 => x"11517080",
  1055 => x"25f43802",
  1056 => x"84050d04",
  1057 => x"02f4050d",
  1058 => x"81ff0bd4",
  1059 => x"0c935380",
  1060 => x"5287fc80",
  1061 => x"c1519ff8",
  1062 => x"2d80c8d4",
  1063 => x"088b3881",
  1064 => x"ff0bd40c",
  1065 => x"8153a1b2",
  1066 => x"04a0eb2d",
  1067 => x"ff135372",
  1068 => x"de387280",
  1069 => x"c8d40c02",
  1070 => x"8c050d04",
  1071 => x"02ec050d",
  1072 => x"810b80cc",
  1073 => x"d00c8454",
  1074 => x"d008708f",
  1075 => x"2a708106",
  1076 => x"51515372",
  1077 => x"f33872d0",
  1078 => x"0ca0eb2d",
  1079 => x"bfe45186",
  1080 => x"b72dd008",
  1081 => x"708f2a70",
  1082 => x"81065151",
  1083 => x"5372f338",
  1084 => x"810bd00c",
  1085 => x"b1538052",
  1086 => x"84d480c0",
  1087 => x"519ff82d",
  1088 => x"80c8d408",
  1089 => x"812e9338",
  1090 => x"72822ebf",
  1091 => x"38ff1353",
  1092 => x"72e438ff",
  1093 => x"145473ff",
  1094 => x"af38a0eb",
  1095 => x"2d83aa52",
  1096 => x"849c80c8",
  1097 => x"519ff82d",
  1098 => x"80c8d408",
  1099 => x"812e0981",
  1100 => x"0693389f",
  1101 => x"a92d80c8",
  1102 => x"d40883ff",
  1103 => x"ff065372",
  1104 => x"83aa2e9e",
  1105 => x"38a1842d",
  1106 => x"a2dd04bf",
  1107 => x"f05186b7",
  1108 => x"2d8053a4",
  1109 => x"b20480c0",
  1110 => x"885186b7",
  1111 => x"2d8054a4",
  1112 => x"830481ff",
  1113 => x"0bd40cb1",
  1114 => x"54a0eb2d",
  1115 => x"8fcf5380",
  1116 => x"5287fc80",
  1117 => x"f7519ff8",
  1118 => x"2d80c8d4",
  1119 => x"085580c8",
  1120 => x"d408812e",
  1121 => x"0981069c",
  1122 => x"3881ff0b",
  1123 => x"d40c820a",
  1124 => x"52849c80",
  1125 => x"e9519ff8",
  1126 => x"2d80c8d4",
  1127 => x"08802e8d",
  1128 => x"38a0eb2d",
  1129 => x"ff135372",
  1130 => x"c638a3f6",
  1131 => x"0481ff0b",
  1132 => x"d40c80c8",
  1133 => x"d4085287",
  1134 => x"fc80fa51",
  1135 => x"9ff82d80",
  1136 => x"c8d408b2",
  1137 => x"3881ff0b",
  1138 => x"d40cd408",
  1139 => x"5381ff0b",
  1140 => x"d40c81ff",
  1141 => x"0bd40c81",
  1142 => x"ff0bd40c",
  1143 => x"81ff0bd4",
  1144 => x"0c72862a",
  1145 => x"70810676",
  1146 => x"56515372",
  1147 => x"963880c8",
  1148 => x"d40854a4",
  1149 => x"83047382",
  1150 => x"2efedb38",
  1151 => x"ff145473",
  1152 => x"fee73873",
  1153 => x"80ccd00c",
  1154 => x"738b3881",
  1155 => x"5287fc80",
  1156 => x"d0519ff8",
  1157 => x"2d81ff0b",
  1158 => x"d40cd008",
  1159 => x"708f2a70",
  1160 => x"81065151",
  1161 => x"5372f338",
  1162 => x"72d00c81",
  1163 => x"ff0bd40c",
  1164 => x"81537280",
  1165 => x"c8d40c02",
  1166 => x"94050d04",
  1167 => x"02e8050d",
  1168 => x"78558056",
  1169 => x"81ff0bd4",
  1170 => x"0cd00870",
  1171 => x"8f2a7081",
  1172 => x"06515153",
  1173 => x"72f33882",
  1174 => x"810bd00c",
  1175 => x"81ff0bd4",
  1176 => x"0c775287",
  1177 => x"fc80d151",
  1178 => x"9ff82d80",
  1179 => x"dbc6df54",
  1180 => x"80c8d408",
  1181 => x"802e8b38",
  1182 => x"80c0a851",
  1183 => x"86b72da5",
  1184 => x"d60481ff",
  1185 => x"0bd40cd4",
  1186 => x"087081ff",
  1187 => x"06515372",
  1188 => x"81fe2e09",
  1189 => x"81069e38",
  1190 => x"80ff539f",
  1191 => x"a92d80c8",
  1192 => x"d4087570",
  1193 => x"8405570c",
  1194 => x"ff135372",
  1195 => x"8025ec38",
  1196 => x"8156a5bb",
  1197 => x"04ff1454",
  1198 => x"73c83881",
  1199 => x"ff0bd40c",
  1200 => x"81ff0bd4",
  1201 => x"0cd00870",
  1202 => x"8f2a7081",
  1203 => x"06515153",
  1204 => x"72f33872",
  1205 => x"d00c7580",
  1206 => x"c8d40c02",
  1207 => x"98050d04",
  1208 => x"02e8050d",
  1209 => x"77797b58",
  1210 => x"55558053",
  1211 => x"727625a3",
  1212 => x"38747081",
  1213 => x"055680f5",
  1214 => x"2d747081",
  1215 => x"055680f5",
  1216 => x"2d525271",
  1217 => x"712e8638",
  1218 => x"8151a695",
  1219 => x"04811353",
  1220 => x"a5ec0480",
  1221 => x"517080c8",
  1222 => x"d40c0298",
  1223 => x"050d0402",
  1224 => x"ec050d76",
  1225 => x"5574802e",
  1226 => x"80c2389a",
  1227 => x"1580e02d",
  1228 => x"51b4b42d",
  1229 => x"80c8d408",
  1230 => x"80c8d408",
  1231 => x"80d3840c",
  1232 => x"80c8d408",
  1233 => x"545480d2",
  1234 => x"e008802e",
  1235 => x"9a389415",
  1236 => x"80e02d51",
  1237 => x"b4b42d80",
  1238 => x"c8d40890",
  1239 => x"2b83fff0",
  1240 => x"0a067075",
  1241 => x"07515372",
  1242 => x"80d3840c",
  1243 => x"80d38408",
  1244 => x"5372802e",
  1245 => x"9d3880d2",
  1246 => x"d808fe14",
  1247 => x"712980d2",
  1248 => x"ec080580",
  1249 => x"d3880c70",
  1250 => x"842b80d2",
  1251 => x"e40c54a7",
  1252 => x"c00480d2",
  1253 => x"f00880d3",
  1254 => x"840c80d2",
  1255 => x"f40880d3",
  1256 => x"880c80d2",
  1257 => x"e008802e",
  1258 => x"8b3880d2",
  1259 => x"d808842b",
  1260 => x"53a7bb04",
  1261 => x"80d2f808",
  1262 => x"842b5372",
  1263 => x"80d2e40c",
  1264 => x"0294050d",
  1265 => x"0402d805",
  1266 => x"0d800b80",
  1267 => x"d2e00c84",
  1268 => x"54a1bc2d",
  1269 => x"80c8d408",
  1270 => x"802e9738",
  1271 => x"80ccd452",
  1272 => x"8051a4bc",
  1273 => x"2d80c8d4",
  1274 => x"08802e86",
  1275 => x"38fe54a7",
  1276 => x"fa04ff14",
  1277 => x"54738024",
  1278 => x"d838738d",
  1279 => x"3880c0b8",
  1280 => x"5186b72d",
  1281 => x"7355adcf",
  1282 => x"04805681",
  1283 => x"0b80d38c",
  1284 => x"0c885380",
  1285 => x"c0cc5280",
  1286 => x"cd8a51a5",
  1287 => x"e02d80c8",
  1288 => x"d408762e",
  1289 => x"09810689",
  1290 => x"3880c8d4",
  1291 => x"0880d38c",
  1292 => x"0c885380",
  1293 => x"c0d85280",
  1294 => x"cda651a5",
  1295 => x"e02d80c8",
  1296 => x"d4088938",
  1297 => x"80c8d408",
  1298 => x"80d38c0c",
  1299 => x"80d38c08",
  1300 => x"802e8181",
  1301 => x"3880d09a",
  1302 => x"0b80f52d",
  1303 => x"80d09b0b",
  1304 => x"80f52d71",
  1305 => x"982b7190",
  1306 => x"2b0780d0",
  1307 => x"9c0b80f5",
  1308 => x"2d70882b",
  1309 => x"720780d0",
  1310 => x"9d0b80f5",
  1311 => x"2d710780",
  1312 => x"d0d20b80",
  1313 => x"f52d80d0",
  1314 => x"d30b80f5",
  1315 => x"2d71882b",
  1316 => x"07535f54",
  1317 => x"525a5657",
  1318 => x"557381ab",
  1319 => x"aa2e0981",
  1320 => x"068e3875",
  1321 => x"51b4832d",
  1322 => x"80c8d408",
  1323 => x"56a9be04",
  1324 => x"7382d4d5",
  1325 => x"2e883880",
  1326 => x"c0e451aa",
  1327 => x"8a0480cc",
  1328 => x"d4527551",
  1329 => x"a4bc2d80",
  1330 => x"c8d40855",
  1331 => x"80c8d408",
  1332 => x"802e83fb",
  1333 => x"38885380",
  1334 => x"c0d85280",
  1335 => x"cda651a5",
  1336 => x"e02d80c8",
  1337 => x"d4088a38",
  1338 => x"810b80d2",
  1339 => x"e00caa90",
  1340 => x"04885380",
  1341 => x"c0cc5280",
  1342 => x"cd8a51a5",
  1343 => x"e02d80c8",
  1344 => x"d408802e",
  1345 => x"8b3880c0",
  1346 => x"f85186b7",
  1347 => x"2daaef04",
  1348 => x"80d0d20b",
  1349 => x"80f52d54",
  1350 => x"7380d52e",
  1351 => x"09810680",
  1352 => x"ce3880d0",
  1353 => x"d30b80f5",
  1354 => x"2d547381",
  1355 => x"aa2e0981",
  1356 => x"06bd3880",
  1357 => x"0b80ccd4",
  1358 => x"0b80f52d",
  1359 => x"56547481",
  1360 => x"e92e8338",
  1361 => x"81547481",
  1362 => x"eb2e8c38",
  1363 => x"80557375",
  1364 => x"2e098106",
  1365 => x"82f93880",
  1366 => x"ccdf0b80",
  1367 => x"f52d5574",
  1368 => x"8e3880cc",
  1369 => x"e00b80f5",
  1370 => x"2d547382",
  1371 => x"2e863880",
  1372 => x"55adcf04",
  1373 => x"80cce10b",
  1374 => x"80f52d70",
  1375 => x"80d2d80c",
  1376 => x"ff0580d2",
  1377 => x"dc0c80cc",
  1378 => x"e20b80f5",
  1379 => x"2d80cce3",
  1380 => x"0b80f52d",
  1381 => x"58760577",
  1382 => x"82802905",
  1383 => x"7080d2e8",
  1384 => x"0c80cce4",
  1385 => x"0b80f52d",
  1386 => x"7080d2fc",
  1387 => x"0c80d2e0",
  1388 => x"08595758",
  1389 => x"76802e81",
  1390 => x"b7388853",
  1391 => x"80c0d852",
  1392 => x"80cda651",
  1393 => x"a5e02d80",
  1394 => x"c8d40882",
  1395 => x"823880d2",
  1396 => x"d8087084",
  1397 => x"2b80d2e4",
  1398 => x"0c7080d2",
  1399 => x"f80c80cc",
  1400 => x"f90b80f5",
  1401 => x"2d80ccf8",
  1402 => x"0b80f52d",
  1403 => x"71828029",
  1404 => x"0580ccfa",
  1405 => x"0b80f52d",
  1406 => x"70848080",
  1407 => x"291280cc",
  1408 => x"fb0b80f5",
  1409 => x"2d708180",
  1410 => x"0a291270",
  1411 => x"80d3800c",
  1412 => x"80d2fc08",
  1413 => x"712980d2",
  1414 => x"e8080570",
  1415 => x"80d2ec0c",
  1416 => x"80cd810b",
  1417 => x"80f52d80",
  1418 => x"cd800b80",
  1419 => x"f52d7182",
  1420 => x"80290580",
  1421 => x"cd820b80",
  1422 => x"f52d7084",
  1423 => x"80802912",
  1424 => x"80cd830b",
  1425 => x"80f52d70",
  1426 => x"982b81f0",
  1427 => x"0a067205",
  1428 => x"7080d2f0",
  1429 => x"0cfe117e",
  1430 => x"29770580",
  1431 => x"d2f40c52",
  1432 => x"59524354",
  1433 => x"5e515259",
  1434 => x"525d5759",
  1435 => x"57adc804",
  1436 => x"80cce60b",
  1437 => x"80f52d80",
  1438 => x"cce50b80",
  1439 => x"f52d7182",
  1440 => x"80290570",
  1441 => x"80d2e40c",
  1442 => x"70a02983",
  1443 => x"ff057089",
  1444 => x"2a7080d2",
  1445 => x"f80c80cc",
  1446 => x"eb0b80f5",
  1447 => x"2d80ccea",
  1448 => x"0b80f52d",
  1449 => x"71828029",
  1450 => x"057080d3",
  1451 => x"800c7b71",
  1452 => x"291e7080",
  1453 => x"d2f40c7d",
  1454 => x"80d2f00c",
  1455 => x"730580d2",
  1456 => x"ec0c555e",
  1457 => x"51515555",
  1458 => x"8051a69f",
  1459 => x"2d815574",
  1460 => x"80c8d40c",
  1461 => x"02a8050d",
  1462 => x"0402ec05",
  1463 => x"0d767087",
  1464 => x"2c7180ff",
  1465 => x"06555654",
  1466 => x"80d2e008",
  1467 => x"8a387388",
  1468 => x"2c7481ff",
  1469 => x"06545580",
  1470 => x"ccd45280",
  1471 => x"d2e80815",
  1472 => x"51a4bc2d",
  1473 => x"80c8d408",
  1474 => x"5480c8d4",
  1475 => x"08802eb8",
  1476 => x"3880d2e0",
  1477 => x"08802e9a",
  1478 => x"38728429",
  1479 => x"80ccd405",
  1480 => x"70085253",
  1481 => x"b4832d80",
  1482 => x"c8d408f0",
  1483 => x"0a0653ae",
  1484 => x"c6047210",
  1485 => x"80ccd405",
  1486 => x"7080e02d",
  1487 => x"5253b4b4",
  1488 => x"2d80c8d4",
  1489 => x"08537254",
  1490 => x"7380c8d4",
  1491 => x"0c029405",
  1492 => x"0d0402e0",
  1493 => x"050d7970",
  1494 => x"842c80d3",
  1495 => x"88080571",
  1496 => x"8f065255",
  1497 => x"53728a38",
  1498 => x"80ccd452",
  1499 => x"7351a4bc",
  1500 => x"2d72a029",
  1501 => x"80ccd405",
  1502 => x"54807480",
  1503 => x"f52d5653",
  1504 => x"74732e83",
  1505 => x"38815374",
  1506 => x"81e52e81",
  1507 => x"f4388170",
  1508 => x"74065458",
  1509 => x"72802e81",
  1510 => x"e8388b14",
  1511 => x"80f52d70",
  1512 => x"832a7906",
  1513 => x"5856769b",
  1514 => x"3880c798",
  1515 => x"08537289",
  1516 => x"387280d0",
  1517 => x"d40b81b7",
  1518 => x"2d7680c7",
  1519 => x"980c7353",
  1520 => x"b1830475",
  1521 => x"8f2e0981",
  1522 => x"0681b638",
  1523 => x"749f068d",
  1524 => x"2980d0c7",
  1525 => x"11515381",
  1526 => x"1480f52d",
  1527 => x"73708105",
  1528 => x"5581b72d",
  1529 => x"831480f5",
  1530 => x"2d737081",
  1531 => x"055581b7",
  1532 => x"2d851480",
  1533 => x"f52d7370",
  1534 => x"81055581",
  1535 => x"b72d8714",
  1536 => x"80f52d73",
  1537 => x"70810555",
  1538 => x"81b72d89",
  1539 => x"1480f52d",
  1540 => x"73708105",
  1541 => x"5581b72d",
  1542 => x"8e1480f5",
  1543 => x"2d737081",
  1544 => x"055581b7",
  1545 => x"2d901480",
  1546 => x"f52d7370",
  1547 => x"81055581",
  1548 => x"b72d9214",
  1549 => x"80f52d73",
  1550 => x"70810555",
  1551 => x"81b72d94",
  1552 => x"1480f52d",
  1553 => x"73708105",
  1554 => x"5581b72d",
  1555 => x"961480f5",
  1556 => x"2d737081",
  1557 => x"055581b7",
  1558 => x"2d981480",
  1559 => x"f52d7370",
  1560 => x"81055581",
  1561 => x"b72d9c14",
  1562 => x"80f52d73",
  1563 => x"70810555",
  1564 => x"81b72d9e",
  1565 => x"1480f52d",
  1566 => x"7381b72d",
  1567 => x"7780c798",
  1568 => x"0c805372",
  1569 => x"80c8d40c",
  1570 => x"02a0050d",
  1571 => x"0402cc05",
  1572 => x"0d7e605e",
  1573 => x"5a800b80",
  1574 => x"d3840880",
  1575 => x"d3880859",
  1576 => x"5c568058",
  1577 => x"80d2e408",
  1578 => x"782e81b8",
  1579 => x"38778f06",
  1580 => x"a0175754",
  1581 => x"73913880",
  1582 => x"ccd45276",
  1583 => x"51811757",
  1584 => x"a4bc2d80",
  1585 => x"ccd45680",
  1586 => x"7680f52d",
  1587 => x"56547474",
  1588 => x"2e833881",
  1589 => x"547481e5",
  1590 => x"2e80fd38",
  1591 => x"81707506",
  1592 => x"555c7380",
  1593 => x"2e80f138",
  1594 => x"8b1680f5",
  1595 => x"2d980659",
  1596 => x"7880e538",
  1597 => x"8b537c52",
  1598 => x"7551a5e0",
  1599 => x"2d80c8d4",
  1600 => x"0880d538",
  1601 => x"9c160851",
  1602 => x"b4832d80",
  1603 => x"c8d40884",
  1604 => x"1b0c9a16",
  1605 => x"80e02d51",
  1606 => x"b4b42d80",
  1607 => x"c8d40880",
  1608 => x"c8d40888",
  1609 => x"1c0c80c8",
  1610 => x"d4085555",
  1611 => x"80d2e008",
  1612 => x"802e9938",
  1613 => x"941680e0",
  1614 => x"2d51b4b4",
  1615 => x"2d80c8d4",
  1616 => x"08902b83",
  1617 => x"fff00a06",
  1618 => x"70165154",
  1619 => x"73881b0c",
  1620 => x"787a0c7b",
  1621 => x"54b3a004",
  1622 => x"81185880",
  1623 => x"d2e40878",
  1624 => x"26feca38",
  1625 => x"80d2e008",
  1626 => x"802eb338",
  1627 => x"7a51add9",
  1628 => x"2d80c8d4",
  1629 => x"0880c8d4",
  1630 => x"0880ffff",
  1631 => x"fff80655",
  1632 => x"5b7380ff",
  1633 => x"fffff82e",
  1634 => x"953880c8",
  1635 => x"d408fe05",
  1636 => x"80d2d808",
  1637 => x"2980d2ec",
  1638 => x"080557b1",
  1639 => x"a2048054",
  1640 => x"7380c8d4",
  1641 => x"0c02b405",
  1642 => x"0d0402f4",
  1643 => x"050d7470",
  1644 => x"08810571",
  1645 => x"0c700880",
  1646 => x"d2dc0806",
  1647 => x"5353718f",
  1648 => x"38881308",
  1649 => x"51add92d",
  1650 => x"80c8d408",
  1651 => x"88140c81",
  1652 => x"0b80c8d4",
  1653 => x"0c028c05",
  1654 => x"0d0402f0",
  1655 => x"050d7588",
  1656 => x"1108fe05",
  1657 => x"80d2d808",
  1658 => x"2980d2ec",
  1659 => x"08117208",
  1660 => x"80d2dc08",
  1661 => x"06057955",
  1662 => x"535454a4",
  1663 => x"bc2d0290",
  1664 => x"050d0402",
  1665 => x"f4050d74",
  1666 => x"70882a83",
  1667 => x"fe800670",
  1668 => x"72982a07",
  1669 => x"72882b87",
  1670 => x"fc808006",
  1671 => x"73982b81",
  1672 => x"f00a0671",
  1673 => x"73070780",
  1674 => x"c8d40c56",
  1675 => x"51535102",
  1676 => x"8c050d04",
  1677 => x"02f8050d",
  1678 => x"028e0580",
  1679 => x"f52d7488",
  1680 => x"2b077083",
  1681 => x"ffff0680",
  1682 => x"c8d40c51",
  1683 => x"0288050d",
  1684 => x"0402f405",
  1685 => x"0d747678",
  1686 => x"53545280",
  1687 => x"71259738",
  1688 => x"72708105",
  1689 => x"5480f52d",
  1690 => x"72708105",
  1691 => x"5481b72d",
  1692 => x"ff115170",
  1693 => x"eb388072",
  1694 => x"81b72d02",
  1695 => x"8c050d04",
  1696 => x"02e8050d",
  1697 => x"77568070",
  1698 => x"56547376",
  1699 => x"24b63880",
  1700 => x"d2e40874",
  1701 => x"2eae3873",
  1702 => x"51aed22d",
  1703 => x"80c8d408",
  1704 => x"80c8d408",
  1705 => x"09810570",
  1706 => x"80c8d408",
  1707 => x"079f2a77",
  1708 => x"05811757",
  1709 => x"57535374",
  1710 => x"76248938",
  1711 => x"80d2e408",
  1712 => x"7426d438",
  1713 => x"7280c8d4",
  1714 => x"0c029805",
  1715 => x"0d0402ec",
  1716 => x"050d80c8",
  1717 => x"d0081751",
  1718 => x"b5802d80",
  1719 => x"c8d40855",
  1720 => x"80c8d408",
  1721 => x"802ea238",
  1722 => x"8b5380c8",
  1723 => x"d4085280",
  1724 => x"d0d451b4",
  1725 => x"d12d80d3",
  1726 => x"90085473",
  1727 => x"802e8a38",
  1728 => x"88155280",
  1729 => x"d0d45173",
  1730 => x"2d029405",
  1731 => x"0d0402dc",
  1732 => x"050d8070",
  1733 => x"5a557480",
  1734 => x"c8d00825",
  1735 => x"b43880d2",
  1736 => x"e408752e",
  1737 => x"ac387851",
  1738 => x"aed22d80",
  1739 => x"c8d40809",
  1740 => x"81057080",
  1741 => x"c8d40807",
  1742 => x"9f2a7605",
  1743 => x"811b5b56",
  1744 => x"547480c8",
  1745 => x"d0082589",
  1746 => x"3880d2e4",
  1747 => x"087926d6",
  1748 => x"38805578",
  1749 => x"80d2e408",
  1750 => x"2781db38",
  1751 => x"7851aed2",
  1752 => x"2d80c8d4",
  1753 => x"08802e81",
  1754 => x"ad3880c8",
  1755 => x"d4088b05",
  1756 => x"80f52d70",
  1757 => x"842a7081",
  1758 => x"06771078",
  1759 => x"842b80d0",
  1760 => x"d40b80f5",
  1761 => x"2d5c5c53",
  1762 => x"51555673",
  1763 => x"802e80cb",
  1764 => x"38741682",
  1765 => x"2bb8da0b",
  1766 => x"80c7a412",
  1767 => x"0c547775",
  1768 => x"311080d3",
  1769 => x"94115556",
  1770 => x"90747081",
  1771 => x"055681b7",
  1772 => x"2da07481",
  1773 => x"b72d7681",
  1774 => x"ff068116",
  1775 => x"58547380",
  1776 => x"2e8a389c",
  1777 => x"5380d0d4",
  1778 => x"52b7d304",
  1779 => x"8b5380c8",
  1780 => x"d4085280",
  1781 => x"d3961651",
  1782 => x"b88e0474",
  1783 => x"16822bb5",
  1784 => x"ce0b80c7",
  1785 => x"a4120c54",
  1786 => x"7681ff06",
  1787 => x"81165854",
  1788 => x"73802e8a",
  1789 => x"389c5380",
  1790 => x"d0d452b8",
  1791 => x"85048b53",
  1792 => x"80c8d408",
  1793 => x"52777531",
  1794 => x"1080d394",
  1795 => x"05517655",
  1796 => x"b4d12db8",
  1797 => x"ab047490",
  1798 => x"29753170",
  1799 => x"1080d394",
  1800 => x"05515480",
  1801 => x"c8d40874",
  1802 => x"81b72d81",
  1803 => x"1959748b",
  1804 => x"24a338b6",
  1805 => x"d3047490",
  1806 => x"29753170",
  1807 => x"1080d394",
  1808 => x"058c7731",
  1809 => x"57515480",
  1810 => x"7481b72d",
  1811 => x"9e14ff16",
  1812 => x"565474f3",
  1813 => x"3802a405",
  1814 => x"0d0402fc",
  1815 => x"050d80c8",
  1816 => x"d0081351",
  1817 => x"b5802d80",
  1818 => x"c8d40880",
  1819 => x"2e893880",
  1820 => x"c8d40851",
  1821 => x"a69f2d80",
  1822 => x"0b80c8d0",
  1823 => x"0cb68e2d",
  1824 => x"90f52d02",
  1825 => x"84050d04",
  1826 => x"02fc050d",
  1827 => x"725170fd",
  1828 => x"2eb03870",
  1829 => x"fd248a38",
  1830 => x"70fc2e80",
  1831 => x"cc38b9f3",
  1832 => x"0470fe2e",
  1833 => x"b73870ff",
  1834 => x"2e098106",
  1835 => x"80c53880",
  1836 => x"c8d00851",
  1837 => x"70802ebb",
  1838 => x"38ff1180",
  1839 => x"c8d00cb9",
  1840 => x"f30480c8",
  1841 => x"d008f405",
  1842 => x"7080c8d0",
  1843 => x"0c517080",
  1844 => x"25a13880",
  1845 => x"0b80c8d0",
  1846 => x"0cb9f304",
  1847 => x"80c8d008",
  1848 => x"810580c8",
  1849 => x"d00cb9f3",
  1850 => x"0480c8d0",
  1851 => x"088c0580",
  1852 => x"c8d00cb6",
  1853 => x"8e2d90f5",
  1854 => x"2d028405",
  1855 => x"0d0402fc",
  1856 => x"050d800b",
  1857 => x"80c8d00c",
  1858 => x"b68e2d8f",
  1859 => x"e32d80c8",
  1860 => x"d40880c8",
  1861 => x"c00c80c7",
  1862 => x"9c519298",
  1863 => x"2d028405",
  1864 => x"0d047180",
  1865 => x"d3900c04",
  1866 => x"00ffffff",
  1867 => x"ff00ffff",
  1868 => x"ffff00ff",
  1869 => x"ffffff00",
  1870 => x"20204368",
  1871 => x"69702d38",
  1872 => x"3a202020",
  1873 => x"20202020",
  1874 => x"50532f32",
  1875 => x"3a000000",
  1876 => x"20203120",
  1877 => x"32203320",
  1878 => x"43202020",
  1879 => x"20202020",
  1880 => x"31203220",
  1881 => x"33203400",
  1882 => x"20203420",
  1883 => x"35203620",
  1884 => x"44202020",
  1885 => x"20202020",
  1886 => x"51205720",
  1887 => x"45205200",
  1888 => x"20203720",
  1889 => x"38203920",
  1890 => x"45202020",
  1891 => x"20202020",
  1892 => x"41205320",
  1893 => x"44204600",
  1894 => x"20204120",
  1895 => x"30204220",
  1896 => x"46202020",
  1897 => x"20202020",
  1898 => x"5a205820",
  1899 => x"43205600",
  1900 => x"3d3d3d20",
  1901 => x"43484950",
  1902 => x"2d382066",
  1903 => x"6f72205a",
  1904 => x"58444f53",
  1905 => x"203d3d3d",
  1906 => x"00000000",
  1907 => x"52657365",
  1908 => x"74000000",
  1909 => x"4c6f6164",
  1910 => x"20526f6d",
  1911 => x"20282e62",
  1912 => x"696e2c20",
  1913 => x"2e636838",
  1914 => x"29201000",
  1915 => x"536f756e",
  1916 => x"64206f6e",
  1917 => x"2f6f6666",
  1918 => x"00000000",
  1919 => x"4b657962",
  1920 => x"6f617264",
  1921 => x"2048656c",
  1922 => x"70000000",
  1923 => x"45786974",
  1924 => x"00000000",
  1925 => x"436c6f63",
  1926 => x"6b205370",
  1927 => x"6565643a",
  1928 => x"20317800",
  1929 => x"436c6f63",
  1930 => x"6b205370",
  1931 => x"6565643a",
  1932 => x"20327800",
  1933 => x"436c6f63",
  1934 => x"6b205370",
  1935 => x"6565643a",
  1936 => x"20337800",
  1937 => x"436c6f63",
  1938 => x"6b205370",
  1939 => x"6565643a",
  1940 => x"20347800",
  1941 => x"3d3d3d20",
  1942 => x"43484950",
  1943 => x"2d382066",
  1944 => x"6f72205a",
  1945 => x"58554e4f",
  1946 => x"203d3d3d",
  1947 => x"00000000",
  1948 => x"524f4d20",
  1949 => x"6c6f6164",
  1950 => x"696e6720",
  1951 => x"6661696c",
  1952 => x"65640000",
  1953 => x"4f4b0000",
  1954 => x"3d3d3d20",
  1955 => x"43484950",
  1956 => x"2d38204b",
  1957 => x"6579626f",
  1958 => x"61726420",
  1959 => x"48454c50",
  1960 => x"203d3d3d",
  1961 => x"00000000",
  1962 => x"3d3d3d3d",
  1963 => x"3d3d3d3d",
  1964 => x"3d3d3d3d",
  1965 => x"3d3d3d3d",
  1966 => x"3d3d3d3d",
  1967 => x"3d3d3d3d",
  1968 => x"3d3d3d3d",
  1969 => x"00000000",
  1970 => x"43686970",
  1971 => x"2d382068",
  1972 => x"61732061",
  1973 => x"20686578",
  1974 => x"206b6579",
  1975 => x"7061642e",
  1976 => x"00000000",
  1977 => x"54686520",
  1978 => x"6d617070",
  1979 => x"696e6720",
  1980 => x"746f2050",
  1981 => x"43206b65",
  1982 => x"79626f61",
  1983 => x"72640000",
  1984 => x"69732066",
  1985 => x"6f6c6c6f",
  1986 => x"77696e67",
  1987 => x"2e000000",
  1988 => x"3d3d3d20",
  1989 => x"43484950",
  1990 => x"2d382043",
  1991 => x"6f726520",
  1992 => x"43726564",
  1993 => x"69747320",
  1994 => x"3d3d3d00",
  1995 => x"43686970",
  1996 => x"2d382063",
  1997 => x"6f726520",
  1998 => x"666f7220",
  1999 => x"5a58554e",
  2000 => x"4f2c2041",
  2001 => x"454f4e2c",
  2002 => x"00000000",
  2003 => x"5a58444f",
  2004 => x"5320616e",
  2005 => x"64205a58",
  2006 => x"444f532b",
  2007 => x"20626f61",
  2008 => x"7264732e",
  2009 => x"00000000",
  2010 => x"4f726967",
  2011 => x"696e616c",
  2012 => x"20636f72",
  2013 => x"65206279",
  2014 => x"3a000000",
  2015 => x"202d2043",
  2016 => x"61727374",
  2017 => x"656e2045",
  2018 => x"6c746f6e",
  2019 => x"20536f72",
  2020 => x"656e7365",
  2021 => x"6e200000",
  2022 => x"506f7274",
  2023 => x"206d6164",
  2024 => x"65206279",
  2025 => x"3a000000",
  2026 => x"202d2041",
  2027 => x"7a65736d",
  2028 => x"626f6700",
  2029 => x"202d2041",
  2030 => x"766c6978",
  2031 => x"41000000",
  2032 => x"496e6974",
  2033 => x"69616c69",
  2034 => x"7a696e67",
  2035 => x"20534420",
  2036 => x"63617264",
  2037 => x"0a000000",
  2038 => x"16200000",
  2039 => x"14200000",
  2040 => x"15200000",
  2041 => x"53442069",
  2042 => x"6e69742e",
  2043 => x"2e2e0a00",
  2044 => x"53442063",
  2045 => x"61726420",
  2046 => x"72657365",
  2047 => x"74206661",
  2048 => x"696c6564",
  2049 => x"210a0000",
  2050 => x"53444843",
  2051 => x"20657272",
  2052 => x"6f72210a",
  2053 => x"00000000",
  2054 => x"57726974",
  2055 => x"65206661",
  2056 => x"696c6564",
  2057 => x"0a000000",
  2058 => x"52656164",
  2059 => x"20666169",
  2060 => x"6c65640a",
  2061 => x"00000000",
  2062 => x"43617264",
  2063 => x"20696e69",
  2064 => x"74206661",
  2065 => x"696c6564",
  2066 => x"0a000000",
  2067 => x"46415431",
  2068 => x"36202020",
  2069 => x"00000000",
  2070 => x"46415433",
  2071 => x"32202020",
  2072 => x"00000000",
  2073 => x"4e6f2070",
  2074 => x"61727469",
  2075 => x"74696f6e",
  2076 => x"20736967",
  2077 => x"0a000000",
  2078 => x"42616420",
  2079 => x"70617274",
  2080 => x"0a000000",
  2081 => x"4261636b",
  2082 => x"00000000",
  2083 => x"00000002",
  2084 => x"00000000",
  2085 => x"00000002",
  2086 => x"00001db0",
  2087 => x"0000039d",
  2088 => x"00000002",
  2089 => x"00001eac",
  2090 => x"0000039d",
  2091 => x"00000002",
  2092 => x"00001dcc",
  2093 => x"00000371",
  2094 => x"00000003",
  2095 => x"00002130",
  2096 => x"00000004",
  2097 => x"00000002",
  2098 => x"00001dd4",
  2099 => x"00001cfe",
  2100 => x"00000001",
  2101 => x"00001dec",
  2102 => x"00000000",
  2103 => x"00000002",
  2104 => x"00001dfc",
  2105 => x"000003b8",
  2106 => x"00000002",
  2107 => x"00001e0c",
  2108 => x"00000800",
  2109 => x"00000002",
  2110 => x"00002480",
  2111 => x"00000000",
  2112 => x"00000002",
  2113 => x"0000249e",
  2114 => x"00000000",
  2115 => x"00000002",
  2116 => x"000024bc",
  2117 => x"00000000",
  2118 => x"00000002",
  2119 => x"000024da",
  2120 => x"00000000",
  2121 => x"00000000",
  2122 => x"00000000",
  2123 => x"00000000",
  2124 => x"00001e14",
  2125 => x"00001e24",
  2126 => x"00001e34",
  2127 => x"00001e44",
  2128 => x"00000002",
  2129 => x"00001e54",
  2130 => x"0000039d",
  2131 => x"00000002",
  2132 => x"00001eac",
  2133 => x"0000039d",
  2134 => x"00000002",
  2135 => x"00001dcc",
  2136 => x"00000371",
  2137 => x"00000003",
  2138 => x"00002130",
  2139 => x"00000004",
  2140 => x"00000002",
  2141 => x"00001dd4",
  2142 => x"00001cfe",
  2143 => x"00000001",
  2144 => x"00001dec",
  2145 => x"00000000",
  2146 => x"00000002",
  2147 => x"00001dfc",
  2148 => x"000003b8",
  2149 => x"00000002",
  2150 => x"00001e0c",
  2151 => x"00000800",
  2152 => x"00000000",
  2153 => x"00000000",
  2154 => x"00000000",
  2155 => x"00000004",
  2156 => x"00001e70",
  2157 => x"000021ac",
  2158 => x"00000004",
  2159 => x"00001e84",
  2160 => x"00002608",
  2161 => x"00000000",
  2162 => x"00000000",
  2163 => x"00000000",
  2164 => x"00000002",
  2165 => x"00001e88",
  2166 => x"0000039c",
  2167 => x"00000002",
  2168 => x"00001ea8",
  2169 => x"0000039c",
  2170 => x"00000002",
  2171 => x"00001ec8",
  2172 => x"0000039c",
  2173 => x"00000002",
  2174 => x"00001ee4",
  2175 => x"0000039c",
  2176 => x"00000002",
  2177 => x"00001f00",
  2178 => x"0000039c",
  2179 => x"00000002",
  2180 => x"00002014",
  2181 => x"0000039c",
  2182 => x"00000002",
  2183 => x"00001d38",
  2184 => x"0000039c",
  2185 => x"00000002",
  2186 => x"00001d50",
  2187 => x"0000039c",
  2188 => x"00000002",
  2189 => x"00001d68",
  2190 => x"0000039c",
  2191 => x"00000002",
  2192 => x"00001d80",
  2193 => x"0000039c",
  2194 => x"00000002",
  2195 => x"00001d98",
  2196 => x"0000039c",
  2197 => x"00000002",
  2198 => x"00002014",
  2199 => x"0000039c",
  2200 => x"00000004",
  2201 => x"00001e84",
  2202 => x"00002608",
  2203 => x"00000000",
  2204 => x"00000000",
  2205 => x"00000000",
  2206 => x"00000002",
  2207 => x"00001f10",
  2208 => x"0000039c",
  2209 => x"00000002",
  2210 => x"00001ea8",
  2211 => x"0000039c",
  2212 => x"00000002",
  2213 => x"00001f2c",
  2214 => x"0000039c",
  2215 => x"00000002",
  2216 => x"00001f4c",
  2217 => x"0000039c",
  2218 => x"00000002",
  2219 => x"00002014",
  2220 => x"0000039c",
  2221 => x"00000002",
  2222 => x"00001f68",
  2223 => x"0000039c",
  2224 => x"00000002",
  2225 => x"00001f7c",
  2226 => x"0000039c",
  2227 => x"00000002",
  2228 => x"00002014",
  2229 => x"0000039c",
  2230 => x"00000002",
  2231 => x"00001f98",
  2232 => x"0000039c",
  2233 => x"00000002",
  2234 => x"00001fa8",
  2235 => x"0000039c",
  2236 => x"00000002",
  2237 => x"00001fb4",
  2238 => x"0000039c",
  2239 => x"00000002",
  2240 => x"00002014",
  2241 => x"0000039c",
  2242 => x"00000004",
  2243 => x"00001e84",
  2244 => x"00002608",
  2245 => x"00000000",
  2246 => x"00000000",
  2247 => x"00000000",
  2248 => x"00000000",
  2249 => x"00000000",
  2250 => x"00000000",
  2251 => x"00000000",
  2252 => x"00000000",
  2253 => x"00000000",
  2254 => x"00000000",
  2255 => x"00000000",
  2256 => x"00000000",
  2257 => x"00000000",
  2258 => x"00000000",
  2259 => x"00000000",
  2260 => x"00000000",
  2261 => x"00000000",
  2262 => x"00000000",
  2263 => x"00000000",
  2264 => x"00000000",
  2265 => x"00000000",
  2266 => x"00000006",
  2267 => x"00000043",
  2268 => x"00000042",
  2269 => x"0000003b",
  2270 => x"0000004b",
  2271 => x"00000033",
  2272 => x"0000001d",
  2273 => x"0000001b",
  2274 => x"0000001c",
  2275 => x"00000023",
  2276 => x"0000002b",
  2277 => x"00000000",
  2278 => x"00000000",
  2279 => x"00000002",
  2280 => x"00002994",
  2281 => x"00001ace",
  2282 => x"00000002",
  2283 => x"000029b2",
  2284 => x"00001ace",
  2285 => x"00000002",
  2286 => x"000029d0",
  2287 => x"00001ace",
  2288 => x"00000002",
  2289 => x"000029ee",
  2290 => x"00001ace",
  2291 => x"00000002",
  2292 => x"00002a0c",
  2293 => x"00001ace",
  2294 => x"00000002",
  2295 => x"00002a2a",
  2296 => x"00001ace",
  2297 => x"00000002",
  2298 => x"00002a48",
  2299 => x"00001ace",
  2300 => x"00000002",
  2301 => x"00002a66",
  2302 => x"00001ace",
  2303 => x"00000002",
  2304 => x"00002a84",
  2305 => x"00001ace",
  2306 => x"00000002",
  2307 => x"00002aa2",
  2308 => x"00001ace",
  2309 => x"00000002",
  2310 => x"00002ac0",
  2311 => x"00001ace",
  2312 => x"00000002",
  2313 => x"00002ade",
  2314 => x"00001ace",
  2315 => x"00000002",
  2316 => x"00002afc",
  2317 => x"00001ace",
  2318 => x"00000004",
  2319 => x"00002084",
  2320 => x"00000000",
  2321 => x"00000000",
  2322 => x"00000000",
  2323 => x"00001c88",
  2324 => x"00000000",
	others => x"00000000"
);

begin

process (clk)
begin
	if (clk'event and clk = '1') then
		if (from_zpu.memAWriteEnable = '1') and (from_zpu.memBWriteEnable = '1') and (from_zpu.memAAddr=from_zpu.memBAddr) and (from_zpu.memAWrite/=from_zpu.memBWrite) then
			report "write collision" severity failure;
		end if;
	
		if (from_zpu.memAWriteEnable = '1') then
			ram(to_integer(unsigned(from_zpu.memAAddr(maxAddrBitBRAM downto 2)))) := from_zpu.memAWrite;
			to_zpu.memARead <= from_zpu.memAWrite;
		else
			to_zpu.memARead <= ram(to_integer(unsigned(from_zpu.memAAddr(maxAddrBitBRAM downto 2))));
		end if;
	end if;
end process;

process (clk)
begin
	if (clk'event and clk = '1') then
		if (from_zpu.memBWriteEnable = '1') then
			ram(to_integer(unsigned(from_zpu.memBAddr(maxAddrBitBRAM downto 2)))) := from_zpu.memBWrite;
			to_zpu.memBRead <= from_zpu.memBWrite;
		else
			to_zpu.memBRead <= ram(to_integer(unsigned(from_zpu.memBAddr(maxAddrBitBRAM downto 2))));
		end if;
	end if;
end process;


end arch;

