12
12
4a
6f
6e
61
73
20
4c
69
6e
64
73
74
65
64
74
00
00
ff
12
8a
64
01
a5
10
6b
00
6c
3b
db
c4
7b
08
3b
80
12
1e
68
3c
a5
08
69
35
d8
96
63
00
43
00
12
3a
a5
0e
d2
32
63
00
8c
40
7c
ff
6b
03
8c
b2
6b
00
4c
00
12
4e
7b
05
7c
ff
12
44
61
00
a4
ee
fb
1e
f0
65
a5
16
f1
1e
f0
55
71
01
7b
01
31
06
12
50
6d
08
6e
05
66
00
6a
01
a5
16
80
d0
d0
e5
70
14
30
6c
12
70
23
44
24
0e
22
f6
23
84
4f
42
12
30
24
46
34
63
12
7a
00
e0
a4
94
6d
28
6e
0a
6c
0a
dd
ea
7d
08
fc
1e
3d
58
12
94
a4
d0
6d
34
6e
19
6c
05
dd
e5
7d
08
fc
1e
3d
4c
12
a6
6d
2d
6e
28
6c
05
dd
e5
7d
08
fc
1e
3d
45
12
b6
a5
15
f0
65
a5
22
f0
33
6c
00
a5
22
fc
1e
f0
65
f0
29
dd
e5
7d
05
7c
01
3c
03
12
ca
6c
0a
ec
9e
12
de
a5
14
60
00
61
00
f1
55
6c
36
00
c1
7c
ff
3c
00
12
ec
12
16
33
00
13
2a
cc
0f
3c
00
13
28
cc
07
7c
01
8c
56
a5
1c
fc
1e
f0
65
40
00
13
28
82
d0
83
e0
73
05
4c
00
13
20
72
14
7c
ff
13
16
a5
0e
d2
32
3f
00
13
38
00
ee
a5
0e
d2
32
73
01
33
3a
13
20
63
00
00
ee
6c
35
8b
30
8b
c5
3f
00
64
63
00
ee
80
40
70
01
80
56
6c
00
a5
1c
fc
1e
f0
55
7c
01
3c
05
13
4c
a5
22
f4
33
23
6c
6c
78
fc
15
fc
07
3c
00
13
62
23
6c
00
ee
a5
23
f0
65
f0
30
6c
37
6b
1b
dc
ba
a5
24
f0
65
f0
30
6c
41
dc
ba
00
ee
46
00
14
00
a5
0e
d5
62
76
ff
46
00
14
00
d5
62
4f
00
14
00
8c
e0
7c
05
8c
65
4f
00
14
02
d5
62
75
fb
66
00
8c
d0
60
00
8b
c0
8b
55
3f
00
13
ba
7c
14
70
01
13
ac
a5
1c
f0
1e
f0
65
70
ff
f0
55
a5
16
40
00
dc
e5
6c
0a
fc
18
a5
14
f0
65
6c
ff
80
c3
f0
55
30
00
13
e4
a5
15
f0
65
70
01
f0
55
6c
00
6b
00
a5
1c
fc
1e
f0
65
30
00
7b
01
7c
01
3c
05
13
e8
3b
00
14
00
74
01
6f
42
00
ee
a5
0e
d2
32
d5
62
63
00
66
00
00
ee
6b
00
6c
03
ec
a1
6b
ff
6c
0c
ec
a1
6b
01
4b
00
14
32
48
01
6b
01
48
78
6b
ff
a5
08
69
35
d8
96
88
b4
d8
96
6c
0a
ec
9e
14
44
36
00
14
44
85
80
66
35
a5
0e
d5
62
00
ee
f0
07
30
00
14
64
60
0a
f0
15
67
00
3d
21
14
5a
6a
ff
14
60
3d
07
14
62
6a
01
67
01
24
66
00
ee
8b
d0
6c
00
89
b0
81
e0
a5
1c
fc
1e
f0
65
40
00
14
82
a5
16
d9
15
89
a4
81
74
d9
15
7c
01
7b
14
3c
05
14
6a
8d
a4
8e
74
4e
30
64
63
00
ee
3c
0c
1e
1e
33
33
3f
61
61
f3
1f
0c
0c
0c
0c
0c
0c
8c
8c
df
07
01
01
01
01
01
01
01
61
e7
e7
83
83
83
83
83
83
83
83
e7
fb
19
01
61
e1
61
01
01
19
fb
9f
86
c6
e6
e6
b6
9e
9e
8e
e6
e4
94
e7
90
f7
87
80
80
80
87
88
88
88
88
af
66
88
48
28
c6
4c
aa
ac
aa
4a
e0
88
c0
88
e0
00
00
18
ff
3c
00
18
3c
ff
81
42
3c
3c
3c
42
3c
5a
5a
7e
7e
00
00
24
3c
24
00
00
18
18
3c
7e
ff
18
18
ff
22
55
88
00
00
00
00
00
00
00
00
00
00
00
00
00
00
00
00
00
00
