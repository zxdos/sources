12
1a
32
2e
30
30
20
43
2e
20
45
67
65
62
65
72
67
20
31
38
2f
38
2d
27
39
31
00
ff
80
03
81
13
a8
e2
f1
55
60
05
a8
e6
f0
55
87
73
86
63
27
86
00
e0
27
a8
6e
40
87
e2
6e
27
87
e1
68
34
69
18
6a
70
6b
00
6c
04
6d
34
27
62
a9
28
da
b8
dc
d8
23
e2
3e
00
12
7e
a8
e6
f0
65
85
00
c4
ff
84
52
25
08
c4
ff
84
52
26
30
60
01
e0
a1
27
f0
36
f7
12
50
8e
60
28
94
6e
64
28
94
27
f0
12
2c
f0
07
40
00
13
22
80
80
80
06
80
06
81
a0
81
06
81
06
80
15
40
00
12
a0
40
01
12
a0
40
ff
12
a0
12
d2
80
90
80
06
80
06
81
b0
81
06
81
06
80
15
40
00
12
bc
40
01
12
bc
40
ff
12
bc
12
d2
a9
28
da
b8
6a
70
6b
00
da
b8
6e
f3
87
e2
6e
04
87
e1
6e
32
28
94
80
80
80
06
80
06
81
c0
81
06
81
06
80
15
40
00
12
ee
40
01
12
ee
40
ff
12
ee
12
56
80
90
80
06
80
06
81
d0
81
06
81
06
80
15
40
00
13
0a
40
01
13
0a
40
ff
13
0a
12
56
a9
28
dc
d8
6c
04
6d
34
dc
d8
6e
cf
87
e2
6e
20
87
e1
6e
19
28
94
12
56
60
3f
28
c2
27
62
a9
28
da
b8
dc
d8
6e
40
87
e3
80
70
80
e2
30
00
12
34
8e
60
28
94
28
a4
00
e0
66
24
67
14
a8
e4
28
00
66
24
67
20
a8
e2
28
00
64
00
65
10
66
01
67
0f
ab
80
d4
60
ab
a0
d5
60
60
03
28
c2
3e
00
13
d8
ab
80
d4
60
ab
a0
d5
60
74
04
75
04
34
60
13
5a
ab
80
d4
60
ab
a0
d5
60
60
03
28
c2
3e
00
13
d8
ab
80
d4
60
ab
a0
d5
60
76
04
36
2d
13
7a
ab
80
d4
60
ab
a0
d5
60
60
03
28
c2
3e
00
13
d8
ab
80
d4
60
ab
a0
d5
60
74
fc
75
fc
34
00
13
98
ab
80
d4
60
ab
a0
d5
60
60
03
28
c2
3e
00
13
d8
ab
80
d4
60
ab
a0
d5
60
76
fc
36
01
13
b8
13
5a
ab
a0
d5
60
ab
c0
d5
60
12
1a
83
70
6e
03
83
e2
84
80
85
90
6e
06
ee
a1
14
44
6e
03
ee
a1
14
5c
6e
08
ee
a1
14
74
6e
07
ee
a1
14
8c
43
03
75
04
43
00
75
fc
43
02
74
04
43
01
74
fc
80
40
81
50
27
d0
82
00
6e
08
80
e2
30
00
14
a4
6e
07
80
20
82
e2
42
05
14
ac
42
06
14
c4
42
07
14
fe
27
62
6e
fc
87
e2
87
31
88
40
89
50
17
62
80
40
81
50
71
04
27
d0
82
00
6e
08
80
e2
30
00
14
04
63
03
75
04
14
20
80
40
81
50
71
fc
27
d0
82
00
6e
08
80
e2
30
00
14
04
63
00
75
fc
14
20
80
40
81
50
70
04
27
d0
82
00
6e
08
80
e2
30
00
14
04
63
02
74
04
14
20
80
40
81
50
70
fc
27
d0
82
00
6e
08
80
e2
30
00
14
04
63
01
74
fc
14
20
27
62
d8
98
8e
f0
00
ee
6e
f0
80
e2
80
31
f0
55
a9
30
d4
58
76
01
61
05
f0
07
40
00
f1
18
14
36
6e
f0
80
e2
80
31
f0
55
a9
38
d4
58
76
04
80
a0
81
b0
27
d0
6e
f0
80
e2
30
00
14
e4
6e
0c
87
e3
80
c0
81
d0
27
d0
6e
f0
80
e2
30
00
14
f6
6e
30
87
e3
60
ff
f0
18
f0
15
14
36
43
01
64
74
43
02
64
00
14
36
82
70
83
70
6e
0c
82
e2
80
a0
81
b0
27
d0
a9
28
6e
f0
80
e2
30
00
15
36
da
b8
42
0c
7b
04
42
00
7b
fc
42
08
7a
04
42
04
7a
fc
da
b8
00
ee
6e
80
f1
07
31
00
15
e6
34
00
15
e6
81
00
83
0e
3f
00
15
68
83
90
83
b5
4f
00
15
9e
33
00
15
86
87
e3
83
80
83
a5
4f
00
15
ce
33
00
15
b6
87
e3
15
e6
83
80
83
a5
4f
00
15
ce
33
00
15
b6
87
e3
83
90
83
b5
4f
00
15
9e
33
00
15
86
87
e3
15
e6
63
40
81
32
41
00
15
e6
da
b8
7b
04
da
b8
6e
f3
87
e2
62
0c
87
21
00
ee
63
10
81
32
41
00
15
e6
da
b8
7b
fc
da
b8
6e
f3
87
e2
62
00
87
21
00
ee
63
20
81
32
41
00
15
e6
da
b8
7a
04
da
b8
6e
f3
87
e2
62
08
87
21
00
ee
63
80
81
32
41
00
15
e6
da
b8
7a
fc
da
b8
6e
f3
87
e2
62
04
87
21
00
ee
c1
f0
80
12
30
00
15
f6
6e
0c
87
e3
82
e3
15
20
da
b8
80
0e
4f
00
16
04
62
04
7a
fc
16
26
80
0e
4f
00
16
10
62
0c
7b
04
16
26
80
0e
4f
00
16
1c
62
08
7a
04
16
26
80
0e
4f
00
15
ee
62
00
7b
fc
da
b8
6e
f3
87
e2
87
21
00
ee
82
70
83
70
6e
30
82
e2
80
c0
81
d0
27
d0
a9
28
6e
f0
80
e2
30
00
16
5e
dc
d8
42
30
7d
04
42
00
7d
fc
42
20
7c
04
42
10
7c
fc
dc
d8
00
ee
6e
80
f1
07
31
00
17
16
34
00
17
16
81
00
83
0e
4f
00
16
90
83
90
83
d5
4f
00
16
c8
33
00
16
ae
87
e3
83
80
83
c5
4f
00
16
fc
33
00
16
e2
87
e3
17
16
83
80
83
c5
4f
00
16
fc
33
00
16
e2
87
e3
83
90
83
d5
4f
00
16
c8
33
00
16
ae
87
e3
17
16
63
40
81
32
41
00
17
16
dc
d8
7d
04
dc
d8
87
e3
6e
cf
87
e2
62
30
87
21
00
ee
63
10
81
32
41
00
17
16
dc
d8
7d
fc
dc
d8
87
e3
6e
cf
87
e2
62
00
87
21
00
ee
63
20
81
32
41
00
17
16
dc
d8
7c
04
dc
d8
87
e3
6e
cf
87
e2
62
20
87
21
00
ee
63
80
81
32
41
00
17
16
dc
d8
7c
fc
dc
d8
87
e3
6e
cf
87
e2
62
10
87
21
00
ee
c1
f0
80
12
30
00
17
28
87
e3
6e
30
87
e3
82
e3
16
48
dc
d8
80
0e
4f
00
17
36
62
90
7c
fc
17
58
80
0e
4f
00
17
42
62
30
7d
04
17
58
80
0e
4f
00
17
4e
62
a0
7c
04
17
58
80
0e
4f
00
17
1e
62
00
7d
fc
dc
d8
6e
4f
87
e2
87
21
00
ee
80
70
6e
03
80
e2
80
0e
81
80
81
94
6e
04
81
e2
41
00
70
01
80
0e
80
0e
80
0e
a8
e8
f0
1e
d8
98
8e
f0
00
ee
6e
00
a9
80
fe
1e
fe
1e
fe
1e
fe
1e
f3
65
ab
e0
fe
1e
fe
1e
fe
1e
fe
1e
f3
55
7e
01
3e
80
17
88
00
ee
82
23
83
33
6e
0f
80
20
81
30
27
d4
80
e2
80
0e
80
0e
a9
40
f0
1e
d2
34
72
04
32
80
17
ae
82
23
73
04
43
40
00
ee
17
ae
70
04
71
04
80
06
80
06
81
06
81
06
81
0e
81
0e
81
0e
81
0e
ab
e0
f1
1e
f1
1e
f0
1e
f0
65
00
ee
a8
e6
f0
65
80
06
f0
55
60
01
e0
a1
17
fa
00
ee
f1
65
6e
01
84
43
82
00
83
10
65
10
83
55
4f
00
82
e5
4f
00
18
26
65
27
82
55
4f
00
18
26
80
20
81
30
84
e4
18
0a
f4
30
d6
7a
76
0c
84
43
82
00
83
10
65
e8
83
55
4f
00
82
e5
4f
00
18
4e
65
03
82
55
4f
00
18
4e
80
20
81
30
84
e4
18
32
f4
30
d6
7a
76
0c
84
43
82
00
83
10
65
64
83
55
4f
00
82
e5
4f
00
18
6e
80
20
81
30
84
e4
18
5a
f4
30
d6
7a
76
0c
84
43
82
00
83
10
65
0a
83
55
4f
00
18
88
81
30
84
e4
18
7a
f4
30
d6
7a
76
0c
f1
30
d6
7a
00
ee
a8
e2
f1
65
81
e4
3f
00
70
01
a8
e2
f1
55
00
ee
a8
e2
f3
65
8e
00
8e
25
4f
00
00
ee
3e
00
18
bc
8e
10
8e
35
4f
00
00
ee
a8
e4
f1
55
00
ee
8e
e3
62
0f
63
ff
61
10
e2
a1
18
de
81
34
31
00
18
ca
61
10
80
34
30
00
18
ca
00
ee
6e
01
00
ee
00
00
00
00
05
00
00
22
63
63
77
7f
3e
1c
00
1c
1e
5d
5d
6f
3e
1c
00
3c
7e
0f
07
0f
7e
3c
00
1c
26
7f
7f
7b
06
1c
00
1e
3f
78
70
78
3f
1e
00
1c
32
7f
7f
6f
30
1c
00
1c
3e
7f
77
63
63
22
00
1c
3e
6f
5d
5d
1e
1c
00
1c
3e
49
77
7f
63
7f
00
00
00
00
08
00
00
00
00
00
00
00
08
08
00
00
00
00
00
00
00
00
00
00
00
00
00
00
00
00
00
00
00
00
00
00
80
00
00
00
80
80
00
00
00
00
00
00
f0
00
00
00
00
00
00
00
80
80
80
80
00
00
00
00
f0
80
80
80
80
80
80
80
f0
00
00
00
80
00
00
00
0c
08
08
08
08
08
08
08
08
08
08
08
08
08
08
0d
0c
08
08
08
08
08
08
08
08
08
08
08
08
08
08
0d
0a
65
05
05
05
05
e5
05
05
e5
05
05
05
05
c5
0a
0a
65
05
05
05
05
e5
05
05
e5
05
05
05
05
c5
0a
0a
05
0c
08
08
0f
05
0c
0d
05
08
08
08
0d
05
0e
0f
05
0c
08
08
0f
05
0c
0d
05
08
08
08
0d
05
0a
0a
05
0a
65
06
05
95
0a
0a
35
05
05
c5
0a
35
05
05
95
0a
65
05
05
95
0a
0a
35
05
06
c5
0a
05
0a
0a
05
0f
05
08
08
08
08
08
0c
08
0f
05
08
08
08
08
08
0f
05
08
08
0c
08
08
08
08
0f
05
0f
05
0a
0a
75
05
b5
05
05
05
05
c5
0a
65
05
b5
05
e5
05
05
e5
05
b5
05
c5
0a
65
05
05
05
05
b5
05
d5
0a
0a
05
0c
08
08
08
08
0d
05
0f
05
0c
08
0f
05
08
0f
05
08
08
0d
05
0f
05
0c
08
08
08
08
0d
05
0a
0f
05
0f
65
05
05
c5
0a
35
e5
95
0a
65
05
b0
05
05
b5
05
c5
0a
35
e5
95
0a
65
05
05
c5
0f
05
0f
07
74
05
d5
08
0f
05
0e
0f
05
08
0f
05
0c
08
08
08
08
0d
05
08
0f
05
08
0f
05
08
0f
75
05
d4
07
0a
05
0a
35
05
05
f5
05
05
b5
05
05
d5
08
08
0d
0c
08
0f
75
05
05
b5
05
05
f5
05
05
95
0a
05
0a
0a
05
08
08
08
0d
05
0c
08
08
08
0d
35
05
c5
0a
0a
65
05
95
0c
08
08
08
0d
05
0c
08
08
0f
05
0a
0a
75
05
06
c5
0a
05
08
08
08
08
08
08
0f
05
08
0f
05
08
08
08
08
08
08
0f
05
0a
65
06
05
d5
0a
0a
05
0c
0d
05
0a
35
05
05
05
05
e5
05
05
f5
05
05
f5
05
05
e5
05
05
05
05
95
0a
05
0c
0d
05
0a
0a
05
08
0f
05
08
08
08
08
08
0f
05
0c
0d
05
08
0f
05
0c
0d
05
08
08
08
08
08
0f
05
08
0f
05
0a
0a
35
05
05
b5
05
05
05
05
05
05
95
0a
0a
35
05
05
95
0a
0a
35
05
05
05
05
05
05
b5
05
05
95
0a
08
08
08
08
08
08
08
08
08
08
08
08
0f
08
08
08
08
08
0f
08
08
08
08
08
08
08
08
08
08
08
08
0f
01
e0
02
10
04
c8
09
e4
0b
f4
0b
b4
09
e5
04
c9
02
13
01
e7
00
07
01
83
03
f0
01
ff
00
ff
00
3f
0f
00
10
80
26
40
4f
20
5f
a0
5d
a0
4f
20
26
40
90
80
cf
00
c0
00
83
00
1f
80
ff
00
fe
00
f8
00
0f
00
1f
80
3f
c0
7f
e0
7f
e0
5f
e0
47
e0
20
c0
90
80
cf
00
c0
80
83
c0
1f
80
ff
00
fe
00
f8
00
