00
e0
cd
7f
ce
7f
8c
d0
8c
e4
a2
a2
6a
00
6b
00
fd
33
f2
65
22
76
a2
88
7a
07
da
b5
a2
a2
7a
08
fe
33
f2
65
22
76
a2
8e
7a
07
da
b4
a2
92
6a
18
6b
08
da
bf
f0
0a
f1
0a
f2
0a
da
bf
6a
15
22
76
a2
a5
f2
55
a2
a2
fc
33
f5
65
83
05
33
00
12
62
84
15
34
00
12
62
85
25
35
00
12
62
66
0c
f6
18
12
6a
6a
15
6b
10
22
76
66
0e
6a
26
6b
08
f6
29
da
b5
f0
0a
12
00
f0
29
da
b5
7a
05
f1
29
da
b5
7a
05
f2
29
da
b5
00
ee
20
20
f8
20
20
00
00
ff
00
ff
ff
ff
03
03
03
ff
ff
c0
c0
c0
c0
c0
00
c0
c0
00
00
00
00
00
00
00
