00
FF
60
01
61
23
62
45
63
67
F3
75
60
00
61
00
62
00
63
00
F3
85
61
04
62
04
22
3C
F3
85
80
10
61
0E
62
04
22
3C
F3
85
80
20
61
18
62
04
22
3C
F3
85
80
30
61
22
62
04
22
3C
00
FD
83
00
83
06
83
06
83
06
83
06
F3
29
D1
25
63
0F
80
32
F0
29
71
05
D1
25
00
EE
