00
ff
6e
0a
00
e0
fe
30
60
04
d0
0a
6d
00
62
04
fe
30
fd
1e
f0
65
61
0f
22
26
72
06
7d
01
3d
0a
12
10
fe
0a
12
04
83
00
83
06
83
06
83
06
83
06
f3
29
d1
25
63
0f
80
32
f0
29
71
05
d1
25
00
ee
