1f
9e
28
63
29
20
41
2e
44
61
75
6d
61
6e
6e
00
e0
00
ff
f2
85
31
aa
00
fd
32
aa
00
fd
ad
d6
f0
55
23
13
23
69
60
00
ad
b5
f0
55
27
6b
ad
b9
60
02
f0
55
27
c9
60
00
ad
cd
f0
55
ad
ce
f0
55
ad
cf
f0
55
ad
d0
f0
55
ad
d1
f0
55
ad
d2
f0
55
ad
d3
f0
55
ad
d4
f0
55
ad
d5
f0
55
27
e7
28
0f
68
08
69
03
24
07
23
c9
60
07
e0
a1
24
55
60
08
e0
a1
24
49
60
0c
e0
a1
24
6f
60
0d
e0
a1
24
63
60
06
e0
a1
24
7d
60
05
e0
a1
24
8d
27
99
ad
b5
f0
65
30
00
12
67
27
d7
ad
b9
f0
65
30
ff
12
a1
12
c1
60
ff
70
01
61
0f
f1
18
61
28
f1
15
f1
07
31
00
12
ad
30
02
12
a3
27
6b
23
c9
24
07
23
c9
12
67
23
c9
28
af
60
ff
70
02
61
0f
f0
18
61
0b
f1
15
f1
07
31
00
12
d1
30
0b
12
c7
ad
d0
f5
65
66
aa
67
aa
f7
75
f0
0a
60
ff
70
01
00
c1
30
40
12
e9
00
fd
ab
44
f5
1e
f0
65
82
00
ab
58
f6
1e
f0
65
83
00
61
06
ab
58
f7
1e
f0
65
a8
ff
f0
1e
d2
36
00
ee
61
ff
71
01
a9
70
f1
1e
f0
65
aa
24
f1
1e
f0
55
31
b3
13
15
00
ee
61
eb
60
ff
70
01
71
01
50
50
13
2d
60
ff
70
01
71
14
50
60
13
37
aa
24
f1
1e
f0
65
87
00
00
ee
61
eb
60
ff
70
01
71
01
50
50
13
4d
60
ff
70
01
71
14
50
60
13
57
aa
24
f1
1e
80
70
f0
55
00
ee
61
fe
67
07
71
02
aa
d8
f1
1e
f0
65
85
00
aa
d9
f1
1e
f0
65
86
00
f1
75
22
f3
f1
85
31
6a
13
6d
00
ee
4a
06
13
a9
4a
07
13
a9
4a
08
13
a9
4a
09
13
a9
4a
0a
13
a9
4a
0b
13
a9
6d
00
87
a0
13
b1
6d
01
87
a0
60
06
87
05
6e
dc
60
ff
7e
24
70
01
50
70
13
b5
00
ee
ab
61
fb
1e
f0
65
8c
00
00
ee
23
bf
61
ff
63
ff
62
ff
73
01
72
01
71
01
3d
00
13
df
ad
ed
13
e1
ae
c5
fe
1e
fc
1e
f1
1e
f0
65
40
ff
13
fd
85
20
85
84
86
30
86
94
87
00
f3
75
22
f3
f3
85
32
02
13
d3
33
02
13
cf
00
ee
61
00
c1
ff
ab
65
f1
1e
f0
65
8a
00
6b
00
23
8b
3a
0b
00
ee
24
29
37
01
00
ee
6a
00
6b
00
23
8b
00
ee
67
00
62
00
61
ff
71
01
aa
24
f1
1e
f0
65
30
06
14
3d
72
01
31
b3
14
2f
32
7e
00
ee
67
01
00
ee
48
11
14
53
23
c9
78
01
23
c9
00
ee
48
00
14
61
23
c9
60
01
88
05
23
c9
00
ee
49
06
14
6d
23
c9
79
01
23
c9
00
ee
49
00
14
7b
23
c9
60
01
89
05
23
c9
00
ee
23
c9
4b
03
14
87
7b
01
14
89
6b
00
23
c9
00
ee
23
bf
61
ff
64
00
63
ff
62
ff
73
01
72
01
71
01
3d
00
14
a5
ad
ed
14
a7
ae
c5
fe
1e
fc
1e
f1
1e
f0
65
40
ff
14
c7
85
20
85
84
86
30
86
94
f3
75
23
29
f3
85
47
06
14
c7
64
01
32
02
14
99
33
02
14
95
34
00
14
d9
4a
0b
15
2b
14
df
4a
0b
15
31
15
2b
60
02
f0
18
23
bf
61
ff
64
00
63
ff
62
ff
73
01
72
01
71
01
3d
00
14
fb
ad
ed
14
fd
ae
c5
fe
1e
fc
1e
f1
1e
f0
65
40
ff
15
19
85
20
85
84
86
30
86
94
f3
75
87
00
23
49
f3
85
32
02
14
ef
33
02
14
eb
25
41
24
07
23
c9
27
6b
00
ee
60
0a
f0
18
00
ee
60
02
f0
18
23
c9
26
81
24
07
23
c9
27
6b
00
ee
61
ff
60
00
71
01
ac
9a
f1
1e
f0
55
ad
18
f1
1e
f0
55
31
7d
15
45
85
80
86
90
75
01
76
01
ac
97
80
50
81
60
f1
55
23
29
ac
8d
f7
1e
f0
65
ac
65
f0
1e
f0
65
82
00
60
00
ac
99
f0
55
32
00
15
c1
00
ee
f3
75
23
29
f3
85
ac
8d
f7
1e
f0
65
ac
79
f0
1e
f1
65
83
00
84
10
52
30
15
af
ac
8d
f7
1e
f0
65
70
01
ac
65
f0
1e
f0
65
82
00
15
c1
52
40
00
ee
ac
8d
f7
1e
f0
65
ac
65
f0
1e
f0
65
82
00
ac
99
f0
65
ac
9a
f0
1e
80
50
f0
55
ac
99
f0
65
ad
18
f0
1e
80
60
f0
55
ac
99
f0
65
70
01
f0
55
60
01
42
01
86
05
42
02
75
01
42
03
76
01
42
04
85
05
ac
97
f1
65
50
50
16
01
51
60
16
01
16
03
15
83
f3
75
23
29
f3
85
ac
8d
f7
1e
f0
65
ac
79
f0
1e
f1
65
83
00
84
10
52
30
16
1f
16
23
52
40
00
ee
26
29
28
37
00
ee
ac
99
f0
65
82
00
60
01
82
05
61
ff
4a
0b
61
00
60
01
f0
18
71
01
ac
9a
f1
1e
f0
65
85
00
ad
18
f1
1e
f0
65
86
00
64
06
f3
75
23
29
80
40
84
70
87
00
23
49
87
40
22
f3
3a
0b
16
6b
67
02
28
69
16
79
ad
d6
f0
65
ad
d7
f0
1e
f0
65
87
00
28
69
f3
85
51
20
16
39
00
ee
61
ff
60
00
71
01
ac
9a
f1
1e
f0
55
ad
18
f1
1e
f0
55
31
7d
16
85
60
00
ac
99
f0
55
ad
96
60
00
f0
55
85
80
86
90
75
01
76
01
ac
97
80
50
81
60
f1
55
f3
75
23
29
f3
85
ad
96
f0
65
81
00
ac
8d
f7
1e
f0
65
80
14
ac
65
f0
1e
f0
65
82
00
32
00
17
13
17
4b
f3
75
23
29
f3
85
ac
8d
f7
1e
f0
65
ac
79
f0
1e
f1
65
83
00
84
10
52
30
17
01
ac
8d
f7
1e
f0
65
70
01
ac
65
f0
1e
f0
65
82
00
17
13
52
40
17
4b
ac
8d
f7
1e
f0
65
ac
65
f0
1e
f0
65
82
00
ac
99
f0
65
40
00
17
2f
ac
9a
f0
1e
80
50
f0
55
ac
99
f0
65
ad
18
f0
1e
80
60
f0
55
ac
99
f0
65
70
01
f0
55
60
01
42
01
86
05
42
02
75
01
42
03
76
01
42
04
85
05
16
d5
ad
96
f0
65
70
01
40
02
17
59
f0
55
16
a3
26
29
00
ee
62
37
ad
97
f7
1e
f0
65
a9
35
d0
25
00
ee
ad
b5
f0
65
81
00
60
01
81
05
60
1e
f0
55
41
1d
17
8b
71
01
87
10
f1
75
27
5d
f1
85
31
1d
17
7d
ad
d6
f0
65
ad
e1
f0
1e
f0
65
f0
15
00
ee
f0
07
30
00
00
ee
ad
b5
f0
65
61
01
80
15
f0
55
87
00
27
5d
ad
d6
f0
65
ad
e1
f0
1e
f0
65
f0
15
00
ee
62
01
ad
b6
f7
1e
f0
65
a9
3a
d2
04
00
ee
67
00
27
bb
67
01
27
bb
67
02
27
bb
00
ee
ad
b9
f0
65
87
00
61
01
80
15
f0
55
27
bb
00
ee
61
ff
64
37
71
01
ad
c4
f1
1e
f0
65
82
00
ad
cd
f1
1e
f0
65
83
00
ad
ba
f3
1e
f0
65
a9
3e
f0
1e
d2
45
31
02
17
eb
00
ee
61
ff
64
37
71
01
ad
c7
f1
1e
f0
65
82
00
ad
d0
f1
1e
f0
65
83
00
ad
ba
f3
1e
f0
65
a9
3e
f0
1e
d2
45
31
05
18
13
00
ee
27
e7
61
03
60
01
81
05
ad
cd
f1
1e
f0
65
40
09
18
4f
70
01
f0
55
18
65
60
00
f0
55
31
00
18
3b
60
00
ad
cd
f0
55
ad
ce
f0
55
ad
cf
f0
55
27
e7
00
ee
28
0f
62
00
72
01
61
06
60
01
81
05
ad
d0
f1
1e
f0
65
40
09
18
85
70
01
f0
55
18
a7
60
00
f0
55
31
00
18
71
60
00
ad
d0
f0
55
ad
d1
f0
55
ad
d2
f0
55
ad
d3
f0
55
ad
d4
f0
55
ad
d5
f0
55
52
70
18
6d
28
0f
00
ee
24
29
37
00
00
ee
6a
0b
63
ff
73
01
62
ff
72
01
85
20
75
01
86
30
76
01
23
29
47
06
18
f5
ad
eb
80
20
f0
55
ad
ec
80
30
f0
55
88
20
89
30
26
81
ad
eb
f0
65
82
00
ad
ec
f0
65
83
00
f3
75
24
29
f3
85
37
00
00
ee
32
11
18
bd
33
06
18
b9
00
ee
7c
fc
c0
c0
cc
cc
f8
fc
0c
0c
cc
cc
cc
cc
c0
c0
fc
7c
cc
cc
0c
0c
fc
f8
cc
cc
cc
cc
cc
cc
fc
fc
00
00
fc
fc
00
00
00
00
00
00
a8
54
a8
54
a8
54
30
78
fc
fc
78
30
c0
c0
c0
c0
c0
60
f0
d0
60
40
a0
a0
a0
40
40
c0
40
40
e0
c0
20
40
80
e0
e0
20
40
20
e0
80
a0
e0
20
20
e0
80
c0
20
e0
60
80
c0
a0
e0
e0
20
40
40
40
e0
a0
40
a0
e0
e0
a0
60
20
c0
07
07
07
07
07
07
07
07
07
07
07
07
07
07
07
07
07
07
07
07
07
06
06
06
06
06
06
06
06
06
06
06
06
06
06
06
06
06
06
07
07
06
06
06
06
06
06
06
06
06
06
06
06
06
06
06
06
06
06
07
07
06
06
06
06
06
06
06
06
06
06
06
06
06
06
06
06
06
06
07
07
06
06
06
06
06
06
06
06
06
06
06
06
06
06
06
06
06
06
07
07
06
06
06
06
06
06
06
06
06
06
06
06
06
06
06
06
06
06
07
07
06
06
06
06
06
06
06
06
06
06
06
06
06
06
06
06
06
06
07
07
06
06
06
06
06
06
06
06
06
06
06
06
06
06
06
06
06
06
07
07
07
07
07
07
07
07
07
07
07
07
07
07
07
07
07
07
07
07
07
07
07
07
07
07
07
07
07
07
07
07
07
07
07
07
07
07
07
07
07
07
06
06
06
06
06
06
06
06
06
06
06
06
06
06
06
06
06
06
07
07
06
06
06
06
06
06
06
06
06
06
06
06
06
06
06
06
06
06
07
07
06
06
06
06
06
06
06
06
06
06
06
06
06
06
06
06
06
06
07
07
06
06
06
06
06
06
06
06
06
06
06
06
06
06
06
06
06
06
07
07
06
06
06
06
06
06
06
06
06
06
06
06
06
06
06
06
06
06
07
07
06
06
06
06
06
06
06
06
06
06
06
06
06
06
06
06
06
06
07
07
06
06
06
06
06
06
06
06
06
06
06
06
06
06
06
06
06
06
07
07
07
07
07
07
07
07
07
07
07
07
07
07
07
07
07
07
07
07
07
00
00
00
01
01
00
00
02
02
00
00
03
03
00
00
04
04
00
00
05
05
00
00
06
06
00
00
07
07
00
00
08
08
00
01
08
09
00
02
08
0a
00
03
08
0b
00
04
08
0c
00
05
08
0d
00
06
08
0e
00
07
08
0f
00
08
08
10
00
09
08
11
00
0a
08
12
00
0b
08
13
00
0c
08
13
01
0d
08
13
02
0e
08
13
03
0f
08
13
04
10
08
13
05
11
08
13
06
12
08
13
07
13
08
06
0c
12
18
1e
24
2a
30
36
3c
42
48
4e
54
5a
60
66
6c
72
78
00
06
0c
12
18
1e
24
2a
30
00
09
12
1b
00
00
00
00
00
00
00
00
00
00
00
00
00
00
00
00
00
00
00
00
00
00
00
00
00
00
00
00
00
00
00
00
00
00
00
00
00
00
00
00
00
00
00
00
00
00
00
00
00
00
00
00
00
00
00
00
00
00
00
01
01
01
01
01
01
01
01
01
01
01
01
01
01
01
01
01
01
01
01
01
01
01
01
01
01
01
01
01
01
01
01
01
01
01
01
01
01
01
01
01
01
01
01
01
01
01
01
01
01
01
01
01
01
01
01
01
01
01
02
02
02
02
02
02
02
02
02
02
02
02
02
02
02
02
02
02
02
02
03
03
03
03
03
03
03
03
03
03
03
03
03
03
03
03
03
03
03
04
04
04
04
04
04
04
04
04
04
04
04
04
04
04
04
04
04
04
05
05
05
05
05
05
05
05
05
05
05
05
05
05
05
05
05
06
06
06
06
06
06
06
06
06
06
06
06
06
06
06
06
06
07
07
07
07
07
07
07
07
07
07
07
07
07
08
08
08
08
08
08
08
08
08
08
08
08
08
09
09
09
09
09
09
09
0a
0a
0a
0a
0a
0a
0a
0b
0b
0b
0b
0b
0b
02
03
04
03
01
02
01
04
01
03
04
02
00
00
00
00
00
00
00
00
04
01
02
01
03
04
03
02
03
01
02
04
00
00
00
00
00
00
00
00
00
02
04
06
08
0a
0c
0e
10
12
00
00
00
00
00
00
00
00
00
00
00
00
00
00
00
00
00
00
00
00
00
00
00
00
00
00
00
00
00
00
00
00
00
00
00
00
00
00
00
00
00
00
00
00
00
00
00
00
00
00
00
00
00
00
00
00
00
00
00
00
00
00
00
00
00
00
00
00
00
00
00
00
00
00
00
00
00
00
00
00
00
00
00
00
00
00
00
00
00
00
00
00
00
00
00
00
00
00
00
00
00
00
00
00
00
00
00
00
00
00
00
00
00
00
00
00
00
00
00
00
00
00
00
00
00
00
00
00
00
00
00
00
00
00
00
00
00
00
00
00
00
00
00
00
00
00
00
00
00
00
00
00
00
00
00
00
00
00
00
00
00
00
00
00
00
00
00
00
00
00
00
00
00
00
00
00
00
00
00
00
00
00
00
00
00
00
00
00
00
00
00
00
00
00
00
00
00
00
00
00
00
00
00
00
00
00
00
00
00
00
00
00
00
00
00
00
00
00
00
00
00
00
00
00
00
00
00
00
00
00
00
00
00
00
00
00
00
00
00
00
00
00
00
00
00
00
00
00
00
00
00
00
00
00
00
00
24
26
28
2a
2c
2e
30
32
34
36
38
3a
3c
3e
40
42
44
46
48
4a
4c
4e
50
52
54
56
58
5a
5c
5e
00
32
2d
28
00
00
05
0a
0f
14
19
1e
23
28
2d
06
0a
0e
67
6b
6f
73
77
7b
00
00
00
00
00
00
00
00
00
00
03
06
09
0c
0f
12
15
18
1b
1e
16
14
12
10
0e
0c
0a
08
06
04
00
00
ff
ff
ff
ff
02
ff
ff
ff
ff
ff
ff
ff
ff
03
ff
ff
ff
ff
ff
ff
ff
ff
01
ff
ff
ff
ff
ff
ff
ff
ff
00
ff
ff
ff
ff
ff
ff
ff
ff
04
ff
ff
ff
ff
ff
ff
ff
ff
05
ff
ff
ff
ff
ff
ff
ff
ff
04
ff
ff
ff
ff
ff
ff
ff
ff
05
ff
ff
ff
ff
ff
04
ff
ff
02
05
ff
ff
ff
ff
04
ff
05
03
ff
ff
ff
ff
ff
ff
ff
05
01
ff
ff
04
ff
ff
ff
ff
ff
00
05
ff
04
ff
ff
ff
ff
00
05
01
04
ff
04
ff
00
05
ff
04
ff
ff
02
05
04
ff
04
02
05
03
ff
ff
ff
05
01
ff
ff
04
ff
05
03
ff
ff
ff
ff
05
05
05
ff
ff
ff
ff
04
ff
ff
04
ff
ff
04
ff
ff
ff
ff
05
05
05
ff
ff
ff
ff
04
ff
ff
04
ff
ff
04
ff
ff
ff
ff
05
05
01
ff
ff
04
ff
00
05
ff
04
ff
ff
04
ff
04
ff
ff
02
05
05
ff
ff
ff
ff
04
ff
ff
04
ff
05
03
ff
ff
ff
ff
00
05
05
04
ff
ff
ff
04
ff
ff
04
ff
ff
02
05
ff
ff
04
05
05
03
ff
ff
ff
05
01
ff
ff
04
ff
ff
04
ff
04
ff
ff
02
01
ff
ff
04
ff
ff
ff
ff
ff
00
05
05
03
ff
04
ff
ff
02
01
ff
ff
04
ff
ff
ff
ff
ff
00
05
05
03
ff
ff
ff
04
ff
00
03
ff
04
ff
05
01
ff
ff
02
05
ff
ff
ff
ff
ff
04
ff
00
03
ff
04
ff
05
01
ff
ff
02
05
ff
ff
ff
04
ff
ff
02
05
01
ff
ff
04
ff
00
05
ff
04
ff
05
03
ff
04
ff
ff
02
05
01
ff
ff
04
ff
00
05
ff
04
ff
05
03
ff
ff
ff
04
00
05
03
04
ff
ff
05
01
ff
ff
04
ff
ff
02
05
ff
ff
04
00
05
03
04
ff
ff
05
01
ff
ff
04
ff
ff
02
05
ff
ff
ff
ff
08
ff
ff
ff
ff
ff
ff
ff
ff
08
ff
ff
ff
ff
ff
ff
ff
ff
08
ff
ff
ff
ff
ff
ff
ff
ff
08
ff
ff
ff
ff
00
00
ff
00
e0
60
0d
61
1b
f0
30
d1
1a
60
00
2f
c4
2f
ce
f1
0a
2f
c4
41
05
1f
e6
41
0c
2f
da
41
0d
2f
e0
2f
c4
1f
ae
f0
30
62
08
63
1b
d2
3a
00
ee
61
10
f1
15
f1
07
31
00
1f
d2
00
ee
30
09
70
01
00
ee
30
00
70
ff
00
ee
00
e0
62
02
f2
18
82
00
60
12
61
0f
a2
00
f1
55
80
20
61
aa
62
aa
f2
75
12
00
