12
16
76
32
2e
30
20
52
61
69
6e
65
73
20
28
63
29
20
31
39
39
31
00
ff
f3
85
8e
20
43
01
12
26
6e
4e
60
00
61
00
a8
6e
f1
55
6c
ff
60
00
61
00
62
00
f2
75
00
e0
60
0b
61
00
62
00
a8
ac
f2
1e
f1
55
72
02
32
78
12
3c
60
00
62
00
a8
64
f2
1e
f1
55
72
02
32
06
12
4c
a8
72
60
26
61
39
63
00
f3
1e
d0
15
63
05
70
08
30
46
12
60
a8
86
60
68
61
02
d0
15
70
08
62
05
f2
1e
d0
15
a8
90
60
68
61
2a
d0
15
70
08
62
05
f2
1e
d0
15
81
e0
81
56
60
64
80
15
a8
1e
f0
33
f2
65
63
5a
64
39
f1
29
d3
45
73
05
f2
29
d3
45
80
e0
a7
bc
f0
55
a7
ce
60
00
61
00
d0
12
70
08
30
60
12
b4
64
02
a7
a4
60
00
d0
4c
a7
b0
60
08
d0
4c
74
0c
34
3e
12
be
67
00
80
70
27
20
77
01
37
05
12
d2
61
32
60
10
a7
de
d0
16
70
08
30
60
12
e2
61
00
60
60
a7
a2
d0
12
71
02
31
38
12
f0
6d
34
24
12
24
1e
24
2c
61
02
a8
16
60
10
d0
18
70
08
30
60
13
06
71
08
31
32
13
04
4c
ff
13
2a
4b
00
63
06
4b
03
63
04
4b
06
63
02
4b
05
63
00
13
38
c3
07
73
01
cc
30
7c
10
8c
34
c3
03
83
5e
a8
5c
f3
1e
f1
65
8b
00
82
10
89
20
80
c0
26
72
26
cc
6a
02
24
3e
67
00
68
00
27
5e
27
80
60
ff
f0
15
60
07
e0
a1
23
aa
60
08
e0
a1
23
c4
60
03
e0
a1
23
de
60
06
e0
a1
23
f8
60
01
e0
a1
23
8c
60
04
e0
a1
23
96
60
0f
e0
a1
6e
02
f0
07
40
00
24
4e
13
5a
60
0f
27
20
80
d0
26
72
00
ee
27
1c
80
d0
26
72
00
ee
80
d0
61
0f
80
12
81
d0
81
05
00
ee
24
12
24
2c
23
9e
70
ff
40
ff
60
00
8d
10
8d
04
24
12
24
2c
60
90
24
36
00
ee
24
12
24
2c
23
9e
70
01
40
0a
60
09
8d
10
8d
04
24
12
24
2c
60
90
24
36
00
ee
24
1e
24
2c
23
9e
71
f0
41
f0
61
00
8d
10
8d
04
24
1e
24
2c
60
90
24
36
00
ee
24
1e
24
2c
23
9e
71
10
41
60
61
50
8d
10
8d
04
24
1e
24
2c
60
90
24
36
00
ee
23
9e
70
60
26
2a
a8
46
d0
14
00
ee
23
9e
80
10
70
0a
26
2a
a8
3e
d0
18
00
ee
80
d0
26
2a
a8
36
d0
18
00
ee
70
ff
30
00
14
36
00
ee
a8
54
fa
1e
f0
65
26
bc
60
6c
61
1c
d0
18
00
ee
24
3e
7a
01
80
90
61
f0
80
12
40
00
14
64
4a
04
14
92
4a
05
15
22
82
a0
3b
00
14
6e
62
08
82
a5
80
b0
80
56
80
56
30
00
14
c0
3b
00
72
ff
80
c0
26
2a
81
24
a8
4a
d0
11
4f
00
15
04
3a
01
15
04
69
00
15
3e
8b
93
60
07
8b
02
80
c0
26
2a
39
16
14
a4
a8
4c
71
04
39
1d
14
ac
a8
4e
71
02
39
15
14
b4
a8
50
71
04
39
1e
14
bc
a8
52
71
02
d0
12
15
22
3b
05
14
d0
63
80
42
08
14
dc
83
56
72
01
14
c6
63
01
42
08
14
dc
83
5e
72
01
14
d2
81
30
80
30
a8
1e
f1
55
a8
1e
80
c0
26
2a
71
03
39
03
14
f6
4a
04
14
f8
3a
05
d0
12
4f
00
15
04
3a
01
15
04
69
00
15
3e
3a
08
15
22
27
5e
60
00
77
01
37
64
15
16
78
01
67
00
70
01
30
03
15
0c
27
5e
6a
00
26
e4
80
e0
81
80
81
74
41
00
70
b0
f0
15
24
3e
00
ee
60
0b
e0
9e
15
34
e0
a1
15
38
00
ee
60
03
f0
18
25
32
00
e0
62
00
63
00
a8
ac
f2
1e
f1
65
72
02
83
14
32
78
15
4a
43
3c
78
01
a8
6e
f1
65
80
74
63
64
80
35
84
f0
34
00
71
01
34
01
70
64
81
84
a8
6e
f1
55
85
00
63
28
64
28
a8
6a
f1
33
f2
65
f0
30
d3
4a
73
0b
f1
30
d3
4a
73
0b
f2
30
d3
4a
a8
6a
f5
33
f2
65
73
0b
f1
30
d3
4a
73
0b
f2
30
d3
4a
27
5e
a7
bc
f0
65
8e
00
4e
02
7e
04
7e
fc
38
00
15
c2
80
56
61
64
81
05
87
15
4f
00
15
cc
25
f6
30
00
12
34
63
01
15
e0
a8
9a
60
2a
61
18
d0
15
70
08
62
05
f2
1e
d0
15
25
f6
63
00
a8
6e
f1
65
82
e0
f3
75
60
0b
e0
a1
15
ea
60
00
e0
a1
15
f0
00
fd
a7
ce
63
02
64
08
d3
48
a7
e6
63
0a
d3
48
a8
a4
63
0e
64
10
d3
47
60
25
24
36
60
0b
e0
a1
16
28
60
00
e0
a1
16
28
d3
47
74
02
44
38
16
06
d3
47
16
0c
00
ee
81
00
6f
f0
81
f2
81
56
6f
0f
80
f2
80
5e
80
5e
80
5e
70
10
71
02
00
ee
70
f0
71
fe
80
56
80
56
80
56
81
5e
80
14
00
ee
a8
ac
81
00
6f
0f
81
f2
81
5e
f1
1e
6f
f0
80
f2
80
56
81
00
81
56
81
56
80
14
80
5e
f0
1e
00
ee
83
00
26
52
f1
65
65
00
30
0b
65
ff
41
00
16
88
61
03
f1
18
16
a4
26
bc
80
30
26
2a
d0
18
80
30
26
52
61
00
80
20
f1
55
80
20
26
bc
80
30
26
2a
d0
18
27
5e
87
54
37
ff
16
b8
48
00
16
b6
78
ff
67
63
16
b8
67
00
27
5e
00
ee
61
0f
80
12
80
5e
80
5e
80
5e
a7
be
f0
1e
00
ee
80
c0
26
52
f1
65
40
0b
15
3e
89
00
80
c0
26
52
80
90
61
01
f1
55
00
ee
63
00
4b
06
63
01
4b
03
63
10
4b
00
63
f0
4b
05
63
ff
81
c0
81
34
6f
f0
81
f2
41
f0
15
3e
41
60
15
3e
81
c0
81
34
6f
0f
81
f2
41
0f
15
3e
41
0a
15
3e
8c
34
26
cc
00
ee
81
a0
17
2a
c1
07
80
56
80
56
40
00
81
56
a8
54
f1
1e
f0
65
85
00
64
03
63
00
a8
64
f3
1e
f0
65
82
00
26
bc
60
04
d0
48
a8
64
f3
1e
80
50
f0
55
26
bc
60
04
d0
48
74
0c
85
20
73
01
33
05
17
36
00
ee
63
69
64
09
a8
6a
f8
33
f2
65
f2
29
d3
45
73
06
a8
6a
f7
33
f2
65
f1
29
d3
45
73
06
f2
29
d3
45
00
ee
80
e0
70
fe
80
56
80
56
61
14
81
05
a8
6a
f1
33
f2
65
f1
30
63
68
64
32
d3
4a
73
0b
f2
30
d3
4a
00
ee
f8
f8
c0
c0
c0
c0
c0
c0
c0
c0
c0
c0
c0
ff
03
03
03
03
03
03
03
03
03
03
03
ff
00
00
00
00
00
00
00
00
00
00
c3
c3
c3
c3
c3
c3
c3
c3
ff
ff
00
00
00
00
ff
ff
c3
c3
00
00
00
00
c3
c3
ff
ff
ff
ff
ff
ff
ff
ff
ff
ff
0f
07
03
03
83
c3
ff
ff
f0
e0
c0
c0
c1
c3
ff
ff
c0
c0
c0
c0
ff
ff
ff
ff
03
03
03
03
ff
ff
c3
c3
c3
c3
c3
c3
ff
ff
ff
ff
c3
c3
c3
c3
c3
c3
00
7e
42
42
42
42
7e
00
00
00
00
00
00
00
00
00
c3
c1
c0
c0
e0
f0
ff
ff
c3
83
03
03
07
0f
ff
ff
00
00
18
3c
3c
18
00
00
00
10
10
70
70
10
10
00
00
18
18
7e
18
00
08
04
04
08
10
20
20
10
1d
15
16
1e
01
02
03
03
06
07
05
08
00
09
03
0a
00
00
00
00
00
00
00
00
00
00
00
00
00
00
a3
a2
e3
a2
aa
bb
92
93
12
3a
bb
a2
b3
22
3a
88
88
88
40
48
d9
92
d2
52
d9
3b
aa
b3
aa
2b
9a
92
9a
91
d9
b4
a4
b4
24
36
ea
aa
ae
a4
e4
ee
8a
ce
89
e9
20
20
70
f8
f8
f8
70
00
0b
00
0b
00
0b
00
0b
00
0b
00
0b
00
0b
00
0b
00
0b
00
0b
00
0b
00
0b
00
0b
00
0b
00
0b
00
0b
00
0b
00
0b
00
0b
00
0b
00
0b
00
0b
00
0b
00
0b
00
0b
00
0b
00
0b
00
0b
00
0b
00
0b
00
0b
00
0b
00
0b
00
0b
00
0b
00
0b
00
0b
00
0b
00
0b
00
0b
00
0b
00
0b
00
0b
00
0b
00
0b
00
0b
00
0b
00
0b
00
0b
00
0b
00
0b
00
0b
00
0b
00
0b
00
0b
00
0b
00
0b
00
0b
00
0b
00
0b
00
