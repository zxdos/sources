00
e0
a2
48
60
00
61
1e
62
00
d2
02
d2
12
72
08
32
40
12
0a
60
00
61
3e
62
02
a2
4a
d0
2e
d1
2e
72
0e
d0
2e
d1
2e
a2
58
60
0b
61
08
d0
1f
70
0a
a2
67
d0
1f
70
0a
a2
76
d0
1f
70
03
a2
85
d0
1f
70
0a
a2
94
d0
1f
12
46
ff
ff
c0
c0
c0
c0
c0
c0
c0
c0
c0
c0
c0
c0
c0
c0
ff
80
80
80
80
80
80
80
80
80
80
80
80
80
ff
81
81
81
81
81
81
81
ff
81
81
81
81
81
81
81
80
80
80
80
80
80
80
80
80
80
80
80
80
80
80
ff
81
81
81
81
81
81
ff
80
80
80
80
80
80
80
ff
81
81
81
81
81
81
ff
81
81
81
81
81
81
ff
ff
